,Unnamed: 0,Name only,page url,Ref count,nb_journal_citations,journalcitation,journal,citation org,citation gov,citation IPCC,citation com,citationipbes,citationguardian,citationautre,org count,gov count,com count,Sci count,IPCC count,percentage of official sources,nbjournaldetected,citationtext_total,Page id,Edit protection,Page lenght (Bytes),DOB,Creator,Total edits,Recent edits,Formated DOB,Year_month,Year
0,0,Medieval cuisine,https://en.wikipedia.org/wiki/Medieval_cuisine,124,3,"['10.1007/s00586-007-0342-x', '10.1484/j.abol.5.102054', '10.2307/2865862', '17390155', None, None, '2200769', None, None]","[['eur spine j'], ['analecta bollandiana'], [' [[speculum ']]",0,0,0,3,0,1,117,0.0,0.0,0.024193548387096774,0.024193548387096774,0.0,0.024193548387096774,3,"['www.nytimes.com', 'books.google.com', 'books.google.com', ['eur spine j'], ['analecta bollandiana'], [' [[speculum ']]",7029997,Allow all users (no expiry set),101475,17 September 2006,Peter Isotalo ,2287,2,2006-09-17,2006-09,2006
1,1,Arab cuisine,https://en.wikipedia.org/wiki/Arab_cuisine,28,0,[],[],1,0,0,16,0,0,11,0.03571428571428571,0.0,0.5714285714285714,0.0,0.0,0.03571428571428571,0,"['books.google.com', 'food.com', 'www.google.com', 'www.nestledessertsarabia.com', 'www.jamaicaobserver.com', 'books.google.com', 'foodspring.com', 'books.google.com', 'mideastfood.about.com', 'www.thestar.com', 'shahiya.com', 'books.google.com', 'www.theglobalist.com', 'www.nytimes.com', 'www.nytimes.com', 'encarta.msn.com', 'nationalfoods.org']",2053043,Allow all users (no expiry set),47418,15 June 2005,128.206.58.214 ,1541,1,2005-06-15,2005-06,2005
2,2,Regional cuisines of medieval Europe,https://en.wikipedia.org/wiki/Regional_cuisines_of_medieval_Europe,19,1,"['10.2307/2598138', None, None]",[['the economic history review']],0,0,0,1,0,0,17,0.0,0.0,0.05263157894736842,0.05263157894736842,0.0,0.05263157894736842,1,"['englishbreakfastsociety.com', ['the economic history review']]",9798488,Allow all users (no expiry set),30834,1 March 2007,Peter Isotalo ,161,0,2007-03-01,2007-03,2007
3,3,European cuisine,https://en.wikipedia.org/wiki/European_cuisine,12,0,[],[],1,0,0,4,0,0,7,0.08333333333333333,0.0,0.3333333333333333,0.0,0.0,0.08333333333333333,0,"['europeword.com', 'books.google.com', 'www.visiteurope.com', 'books.google.com', 'www.lordsandladies.org']",524762,Allow all users (no expiry set),26333,13 March 2004,Mkweise ,1695,21,2004-03-13,2004-03,2004
4,4,List of cuisines,https://en.wikipedia.org/wiki/List_of_cuisines,4,0,[],[],0,0,0,3,0,0,1,0.0,0.0,0.75,0.0,0.0,0.0,0,"['oxforddictionaries.com', 'thefreedictionary.com', 'www.merriam-webster.com']",265366,Allow all users (no expiry set),24388,11 July 2003,142.177.97.12 ,1156,2,2003-07-11,2003-07,2003
5,5,Byzantine cuisine,https://en.wikipedia.org/wiki/Byzantine_cuisine,6,1,"['10.1017/s1380203800001756', None, None]",[['archaeological dialogues ']],0,0,0,3,0,0,2,0.0,0.0,0.5,0.16666666666666666,0.0,0.16666666666666666,1,"['books.google.com', 'books.google.com', 'www.reuters.com', ['archaeological dialogues ']]",5771126,Allow all users (no expiry set),9780,30 June 2006,NickOfCyprus ,192,0,2006-06-30,2006-06,2006
6,6,French cuisine,https://en.wikipedia.org/wiki/French_cuisine,38,1,"['10.2307/1843902', None, None]",[['the american historical review']],3,0,0,9,0,1,24,0.07894736842105263,0.0,0.23684210526315788,0.02631578947368421,0.0,0.10526315789473684,1,"['www.frenchentree.com', 'www.bibliotheque-dauphinoise.com', 'travelfoodatlas.com', 'cheznoscousins.com', 'www.leershistorique.com', 'www.nice-cooking.com', 'www.dallasnews.com', 'french-country-decor-guide.com', 'www.joyeux-noel.com', 'www.unesco.org', 'www.ambafrance-at.org', 'menus.nypl.org', ['the american historical review']]",11002,Allow all users (no expiry set),80853,22 August 2001,47.83.107.xxx ,4451,2,2001-08-22,2001-08,2001
7,7,Catalan cuisine,https://en.wikipedia.org/wiki/Catalan_cuisine,25,1,"['10.2752/175174409x456737', None, None]",[[' food']],0,0,0,11,0,0,13,0.0,0.0,0.44,0.04,0.0,0.04,1,"['www.llibreriaona.com', 'www.catalannews.com', 'books.google.com', 'books.google.com', 'www.comunitatvalenciana.com', 'books.google.com', 'www.comunitatvalenciana.com', 'www.google.com', 'www.catalannews.com', 'articles.economictimes.indiatimes.com', 'www.nytimes.com', [' food']]",71058,Allow all users (no expiry set),22354,13 August 2002,Perique des Palottes ,447,1,2002-08-13,2002-08,2002
8,8,Early modern European cuisine,https://en.wikipedia.org/wiki/Early_modern_European_cuisine,20,1,"['10.1353/jwh.2016.0020', None, None]",[['journal of world history']],0,0,0,1,0,0,18,0.0,0.0,0.05,0.05,0.0,0.05,1,"['www.houseofbols.com', ['journal of world history']]",10928780,Allow all users (no expiry set),23939,27 April 2007,Peter Isotalo ,206,3,2007-04-27,2007-04,2007
9,9,List of historical cuisines,https://en.wikipedia.org/wiki/List_of_historical_cuisines,2,0,[],[],0,0,0,1,0,0,1,0.0,0.0,0.5,0.0,0.0,0.0,0,['docs.google.com'],44796268,Allow all users (no expiry set),2041,21 December 2014,Chiswick Chap ,32,0,2014-12-21,2014-12,2014
10,10,Mughlai cuisine,https://en.wikipedia.org/wiki/Mughlai_cuisine,8,1,"['10.7208/chicago/9780226243276.003.0004', None, None]",[['university of chicago press']],0,0,0,6,0,0,1,0.0,0.0,0.75,0.125,0.0,0.125,1,"['www.telegraphindia.com', 'gulfnews.com', 'www.dawn.com', 'www.outlookindia.com', 'www.indiatimes.com', 'www.thebetterindia.com', ['university of chicago press']]",13107093,Allow all users (no expiry set),9857,5 September 2007,Randhirreddy ,472,1,2007-09-05,2007-09,2007
11,11,Sicilian cuisine,https://en.wikipedia.org/wiki/Sicilian_cuisine,17,0,[],[],0,0,0,5,0,0,12,0.0,0.0,0.29411764705882354,0.0,0.0,0.0,0,"['www.etnasicilytouring.com', 'books.google.com', 'books.google.com', 'www.mangiabedda.com', 'www.tesorichicago.com']",44808,Allow all users (no expiry set),14208,18 March 2002,Zisa ,322,0,2002-03-18,2002-03,2002
12,12,Haute cuisine,https://en.wikipedia.org/wiki/Haute_cuisine,6,0,[],[],0,0,0,1,0,0,5,0.0,0.0,0.16666666666666666,0.0,0.0,0.0,0,['books.google.com'],334079,Allow all users (no expiry set),8411,3 October 2003,UninvitedCompany ,316,0,2003-10-03,2003-10,2003
13,13,Roman cuisine,https://en.wikipedia.org/wiki/Roman_cuisine,17,0,[],[],0,0,0,1,0,0,16,0.0,0.0,0.058823529411764705,0.0,0.0,0.0,0,['sweets.seriouseats.com'],25882073,Allow all users (no expiry set),9569,20 January 2010,Theologiae ,347,0,2010-01-20,2010-01,2010
14,14,Italian cuisine,https://en.wikipedia.org/wiki/Italian_cuisine,235,0,[],[],5,2,0,92,0,3,133,0.02127659574468085,0.00851063829787234,0.39148936170212767,0.0,0.0,0.029787234042553193,0,"['www.uibm.gov', 'nla.gov', 'www.webfoodculture.com', 'educalingo.com', 'www.theatlantic.com', 'www.unionalimentari.com', 'books.google.com', 'books.google.com', 'www.thrillist.com', 'it.yougov.com', 'tasteatlas.com', 'tableagent.com', 'www.americanheritage.com', 'britannica.com', 'rusticocooking.com', 'www.fondazioneslowfood.com', 'notitarde.com', 'www.delallo.com', 'it.healthy-food-near-me.com', 'yourguidetoitaly.com', 'winefolly.com', 'books.google.com', 'educalingo.com', 'www.fondazioneslowfood.com', 'italianfood.about.com', 'lacucinaitaliana.com', 'www.slowfood.com', 'www.aspenbusinessjournal.com', 'sweets.seriouseats.com', 'www.americanheritage.com', 'www.lomejordelagastronomia.com', 'www.delallo.com', 'thestreet.com', 'www.moldrek.com', 'www.slowfood.com', 'toscanaslc.com', 'www.annamariavolpi.com', 'www.greatitalianchefs.com', 'books.google.com', 'it.yougov.com', 'books.google.com', 'books.google.com', 'www.italianfoodexcellence.com', 'books.google.com', 'blog.tuscany-cooking-class.com', 'blog.tuscany-cooking-class.com', 'italianowine.com', 'books.google.com', 'sallybernstein.com', 'www.ristonews.com', 'eritrealive.com', 'giornalevinocibo.com', 'thestreet.com', 'books.google.com', 'it.ripleybelieves.com', 'www.epicurean.com', 'hillmanwonders.com', 'www.forbes.com', 'www.lifeinitaly.com', 'books.google.com', 'yosoymukenio.blogspot.com', 'www.thejakartapost.com', 'magazine.luxuryretreats.com', 'knopfdoubleday.com', 'edition.cnn.com', 'books.google.com', 'www.silviocicchi.com', 'tasteatlas.com', 'it.encyclopedia-titanica.com', 'www.alfemminile.com', 'www.lifeinitaly.com', 'www.oliveoiltimes.com', 'www.nytimes.com', 'www.deliciousitaly.com', 'books.google.com', 'fresco.irinox.com', 'www.deliciousitaly.com', 'winefolly.com', 'www.indigoguide.com', 'www.italianfoodexcellence.com', 'www.chowhound.com', 'www.eataly.com', 'www.hotelposeidontortoreto.com', 'www.nytimes.com', 'www.baristabasics.com', 'books.google.com', 'magazine.luxuryretreats.com', 'www.malta-turismo.com', 'books.google.com', 'www.apreroma.com', 'greatitalianchefs.com', 'books.google.com', 'www.timescolonist.com', 'www.bbcgoodfood.com', 'www.inta.org', 'r0.unctad.org', 'www.pizzanapoletana.org', 'www.genteditalia.org', 'expo2015.org']",3735620,Allow all users (no expiry set),152002,16 January 2006,AKeen ,4829,22,2006-01-16,2006-01,2006
15,15,Bavarian cuisine,https://en.wikipedia.org/wiki/Bavarian_cuisine,9,0,[],[],0,0,0,3,0,0,6,0.0,0.0,0.3333333333333333,0.0,0.0,0.0,0,"['books.google.com', 'books.google.com', 'www.nytimes.com']",22946736,Allow all users (no expiry set),13145,25 May 2009,Pitoutom ,165,0,2009-05-25,2009-05,2009
16,16,Hyderabadi cuisine,https://en.wikipedia.org/wiki/Hyderabadi_cuisine,29,0,[],[],0,0,0,26,0,0,3,0.0,0.0,0.896551724137931,0.0,0.0,0.0,0,"['books.google.com', 'www.thehindu.com', 'articles.timesofindia.indiatimes.com', 'www.slate.com', 'www.newindianexpress.com', 'www.thehindu.com', 'www.deccanchronicle.com', 'www.thehindu.com', 'books.google.com', 'recipes.timesofindia.com', 'www.thenewsminute.com', 'yummyindiankitchen.com', 'books.google.com', 'khanapakana.com', 'www.newindianexpress.com', 'www.deccanchronicle.com', 'www.nytimes.com', 'timesofindia.indiatimes.com', 'food.ndtv.com', 'www.deccanchronicle.com', 'india.blogs.nytimes.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'books.google.com', 'www.newindianexpress.com', 'www.rediff.com']",11659590,Allow all users (no expiry set),19736,8 June 2007,Randhirreddy ,650,4,2007-06-08,2007-06,2007
17,17,Cuisine,https://en.wikipedia.org/wiki/Cuisine,15,0,[],[],1,0,0,8,0,1,5,0.06666666666666667,0.0,0.5333333333333333,0.0,0.0,0.06666666666666667,0,"['www.britannica.com', 'books.google.com', 'www.kraft.com', 'www.chinadaily.com', 'www.merriam-webster.com', 'www.scienceofcooking.com', 'query.nytimes.com', 'www.ricearoni.com', 'web-japan.org']",6656,Allow all users (no expiry set),20724,26 October 2001,202.36.170.xxx ,1212,3,2001-10-26,2001-10,2001
18,18,Sichuan cuisine,https://en.wikipedia.org/wiki/Sichuan_cuisine,15,1,"['10.1016/j.fshw.2019.03.008', None, None]",[['food science and human wellness ']],1,0,0,7,0,0,6,0.06666666666666667,0.0,0.4666666666666667,0.06666666666666667,0.0,0.13333333333333333,1,"['mychinesesoulfood.com', 'www.britannica.com', 'www.flavorandfortune.com', 'blogs.wsj.com', 'www.phaidon.com', 'www.aboluowang.com', 'www.chinasichuanfood.com', 'unesdoc.unesco.org', ['food science and human wellness ']]",27908,Allow all users (no expiry set),19143,5 November 2001,24.4.254.xxx ,661,47,2001-11-05,2001-11,2001
19,19,Mediterranean cuisine,https://en.wikipedia.org/wiki/Mediterranean_cuisine,91,13,"['10.1016/j.dib.2017.05.007', '10.1093/ajcn/61.6.1313s', '10.1024/0300-9831.71.3.141', '10.1016/j.tig.2006.07.008', '10.1007/bf02904806', '10.21273/hortsci.42.5.1093', '10.1093/ajcn/61.6.1402s', '10.1093/aob/mcp298', '10.1126/science.1124635', '10.1016/j.appet.2018.10.022', '10.13140/rg.2.1.2690.8327', '10.1007/bf00029633', '10.1080/07409710.2017.1270646', '28560272', '7754981', '11582834', '16872714', None, None, '7754995', '20034966', '16574859', None, None, None, None, '5435575', None, None, None, None, None, None, '2826248', None, None, None, None, None]","[['data in brief '], ['american journal of clinical nutrition '], ['int j vitam nutr res '], ['trends in genetics '], ['economic botany '], ['hortscience '], ['american journal of clinical nutrition '], ['ann bot '], ['science '], ['appetite '], ['universidad de córdoba '], ['euphytica '], ['food and foodways ']]",6,0,0,24,0,2,46,0.06593406593406594,0.0,0.26373626373626374,0.14285714285714285,0.0,0.2087912087912088,13,"['books.google.com', 'www.visitportugal.com', 'books.google.com', 'books.google.com', 'www.theatlantic.com', 'books.google.com', 'books.google.com', 'tableagent.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'play.google.com', 'www.latimes.com', 'books.google.com', 'books.google.com', 'www.ft.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'tasteporto.com', 'books.google.com', 'food.com', 'www.spanish-food.org', 'www.iemed.org', 'www.fao.org', 'faostat.fao.org', 'www.cabdirect.org', 'www.diabetes.org', ['data in brief '], ['american journal of clinical nutrition '], ['int j vitam nutr res '], ['trends in genetics '], ['economic botany '], ['hortscience '], ['american journal of clinical nutrition '], ['ann bot '], ['science '], ['appetite '], ['universidad de córdoba '], ['euphytica '], ['food and foodways ']]",1342098,Allow all users (no expiry set),56847,29 December 2004,62.74.2.11 ,1159,5,2004-12-29,2004-12,2004
20,20,Cuisine of Abruzzo,https://en.wikipedia.org/wiki/Cuisine_of_Abruzzo,28,0,[],[],1,0,0,19,0,0,8,0.03571428571428571,0.0,0.6785714285714286,0.0,0.0,0.03571428571428571,0,"['articles.philly.com', 'books.google.com', 'articles.philly.com', 'www.hotelposeidontortoreto.com', 'books.google.com', 'italy.com', 'www.delallo.com', 'www.bompensaoliveoil.com', 'www.lifeinabruzzo.com', 'www.academiabarilla.com', 'books.google.com', 'www.delallo.com', 'books.google.com', 'www.ashbytreats.com', 'lifeinabruzzo.com', 'books.google.com', 'issuu.com', 'www.huffingtonpost.com', 'www.cookaround.com', 'abruzzomoliseheritagesociety.org']",43385749,Allow all users (no expiry set),23383,24 July 2014,Pete Maverick ,165,1,2014-07-24,2014-07,2014
21,21,Balkan cuisine,https://en.wikipedia.org/wiki/Balkan_cuisine,18,1,"['10.2307/628548', None, None]",[['the journal of hellenic studies ']],1,0,0,14,0,0,2,0.05555555555555555,0.0,0.7777777777777778,0.05555555555555555,0.0,0.1111111111111111,1,"['books.google.com', 'books.google.com', 'theculturetrip.com', 'www.washingtonpost.com', 'balkaninsight.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.npr.org', ['the journal of hellenic studies ']]",49733604,Allow all users (no expiry set),10844,11 March 2016,Polly Tunnel ,82,5,2016-03-11,2016-03,2016
22,22,List of European cuisines,https://en.wikipedia.org/wiki/List_of_European_cuisines,29,0,[],[],2,1,0,19,0,1,6,0.06896551724137931,0.034482758620689655,0.6551724137931034,0.0,0.0,0.10344827586206896,0,"['www.cia.gov', 'thefreedictionary.com', 'ukraine.com', 'sallybernstein.com', 'ultimate-guide-to-greek-food.com', 'homecooking.about.com', 'food-links.com', 'indigoguide.com', 'britannica.com', 'europeword.com', 'cooking-advices.com', 'buzzle.com', 'www.dallasnews.com', 'www.colonialvoyage.com', 'books.google.com', 'french-country-decor-guide.com', 'books.google.com', 'goeasteurope.about.com', 'ukrainetrek.com', 'rusticocooking.com', 'www.unesco.org', 'www.cac-biodiversity.org']",39488476,Allow all users (no expiry set),31775,26 May 2013,The Transhumanist ,311,7,2013-05-26,2013-05,2013
23,23,Chinese cuisine,https://en.wikipedia.org/wiki/Chinese_cuisine,70,7,"['10.1038/514s58a', '10.1016/j.jef.2015.11.004', '10.1038/s41477-018-0141-x', '10.1080/10942912.2017.1382507', '10.1016/s0168-1605(00)00523-7', '10.17730/humo.45.2.4034u85x3058m025', '10.1016/j.jef.2016.08.003', '25368889', None, '29725102', None, '11322691', None, None, None, None, None, None, None, None, None]","[['nature'], ['journal of ethnic foods'], ['nature plants'], ['international journal of food properties '], ['international journal of food microbiology'], ['human organization '], ['journal of ethnic foods']]",5,0,0,29,0,0,29,0.07142857142857142,0.0,0.4142857142857143,0.1,0.0,0.17142857142857143,7,"['simplechinesefood.com', 'www.theatlantic.com', 'chinesefood.about.com', 'books.google.com', 'www.eatingchina.com', 'www.chinatoday.com', 'books.google.com', 'www.sciencedaily.com', 'languageoffood.blogspot.com', 'wayoftheeating.wordpress.com', 'www.flavorandfortune.com', 'books.google.com', 'kaleidoscope.cultural-china.com', 'books.google.com', 'books.google.com', 'supchina.com', 'beautyfujian.com', 'www.economist.com', 'www.yumofchina.com', 'www.nytimes.com', 's.visitbeijing.com', 'books.google.com', 'books.google.com', 'www.dummies.com', 'www.flavorandfortune.com', 'wayoftheeating.wordpress.com', 'data.eastmoney.com', 'books.google.com', 'www.geog.com', 'www.worldcat.org', 'www.ibiblio.org', 'dictionary.cambridge.org', 'ethnomed.org', 'www.ibiblio.org', ['nature'], ['journal of ethnic foods'], ['nature plants'], ['international journal of food properties '], ['international journal of food microbiology'], ['human organization '], ['journal of ethnic foods']]",6583,Allow all users (no expiry set),58674,25 September 2001,Dmerrill ,5240,10,2001-09-25,2001-09,2001
24,24,Spanish cuisine,https://en.wikipedia.org/wiki/Spanish_cuisine,83,8,"['10.5944/etfiii.16.2003.3689', '10.1080/14636204.2013.916027', '10.30687/978-88-6969-302-1/006', '10.3989/chdj.2017.019', '10.3390/nu10091234', '10.1057/9781137324054', '10.7827/turkishstudies.12900', None, None, None, None, '30189597', None, None, None, None, None, None, '6164545', None, None]","[['[[universidad nacional de educación a distancia', 'espacio'], ['journal of spanish cultural studies', '[[routledge'], ['edizioni ca'], ['culture '], ['nutrients'], ['[[palgrave macmillan'], ['turkish studies']]",2,0,0,34,0,1,38,0.024096385542168676,0.0,0.40963855421686746,0.0963855421686747,0.0,0.12048192771084337,7,"['books.google.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'www.korespa.com', 'elpais.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.elespanol.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'theculturetrip.com', 'www.josemadeinspain.com', 'www.latimes.com', 'books.google.com', 'www.saveur.com', 'diariodegastronomia.com', 'www.elespanol.com', 'academiaaragonesadegastronomia.com', 'books.google.com', 'clic-books.com', 'www.nytimes.com', 'www.revistagq.com', 'www.foodandwine.com', 'elcomidista.elpais.com', 'books.google.com', 'books.google.com', 'www.revistadelibros.com', 'elcomidista.elpais.com', 'www.latimes.com', 'www.spanish-food.org', 'www.eurofir.org', ['[[universidad nacional de educación a distancia', 'espacio'], ['journal of spanish cultural studies', '[[routledge'], ['edizioni ca'], ['culture '], ['nutrients'], ['[[palgrave macmillan'], ['turkish studies']]",27669,Allow all users (no expiry set),64541,22 September 2001,137.110.9.xxx ,2419,0,2001-09-22,2001-09,2001
25,25,Arbëreshë cuisine,https://en.wikipedia.org/wiki/Arb%C3%ABresh%C3%AB_cuisine,1,0,[],[],0,0,0,1,0,0,0,0.0,0.0,1.0,0.0,0.0,0.0,0,['books.google.com'],56594785,Allow all users (no expiry set),1118,15 February 2018,Iaof2017 ,14,0,2018-02-15,2018-02,2018
26,26,Venetian cuisine,https://en.wikipedia.org/wiki/Venetian_cuisine,2,0,[],[],0,0,0,0,0,0,2,0.0,0.0,0.0,0.0,0.0,0.0,0,[],26348119,Allow all users (no expiry set),14491,26 February 2010,Theologiae ,150,0,2010-02-26,2010-02,2010
27,27,Indian cuisine,https://en.wikipedia.org/wiki/Indian_cuisine,266,1,"['10.1016/j.yclnex.2019.05.004', None, None]",[['clinical nutrition experimental ']],6,2,0,208,0,2,47,0.022556390977443608,0.007518796992481203,0.7819548872180451,0.0037593984962406013,0.0,0.03383458646616541,1,"['www.food.gov', 'www.food.gov', 'hebbarskitchen.com', 'www.tribuneindia.com', 'www.onmanorama.com', 'www.thehindu.com', 'books.google.com', 'medium.com', 'books.google.com', 'www.bestindianfoodcatering.com', 'www.archanaskitchen.com', 'www.cookwithmanali.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'vice.com', 'hebbarskitchen.com', 'books.google.com', 'books.google.com', 'www.telegraphindia.com', 'books.google.com', 'books.google.com', 'www.archanaskitchen.com', 'books.google.com', 'books.google.com', 'articles.economictimes.indiatimes.com', 'www.mygingergarlickitchen.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'theflavoursofhistory.com', 'lulu.com', 'indiasite.com', 'hoggngulp.blogspot.com', 'books.google.com', 'books.google.com', 'recipes.timesofindia.com', 'india9.com', 'books.google.com', 'www.enhanceyourpalate.com', 'www.archanaskitchen.com', 'm.recipes.timesofindia.com', 'indianfoodforever.com', 'rediff.com', 'books.google.com', 'business.google.com', 'articles.timesofindia.indiatimes.com', 'books.google.com', 'konkanifoodrecipes.com', 'indianexpress.com', 'm.recipes.timesofindia.com', 'books.google.com', 'mapsofindia.com', 'www.archanaskitchen.com', 'www.archanaskitchen.com', 'food-india.com', 'books.google.com', 'books.google.com', 'books.google.com', 'articles.timesofindia.indiatimes.com', 'bhavnaskitchen.com', 'www.temptingtreat.com', 'traveller.outlookindia.com', 'books.google.com', 'books.google.com', 'kalimirchbysmita.com', '10keythings.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.vegrecipesofindia.com', 'www.foodvedam.com', 'www.archanaskitchen.com', 'myvegetarianroots.com', 'www.business-standard.com', 'books.google.com', 'www.archanaskitchen.com', 'books.google.com', 'maayeka.com', 'books.google.com', 'foodtourindelhi.com', 'www.hindu.com', 'recipes.timesofindia.com', 'www.newindianexpress.com', 'www.archanaskitchen.com', 'ministryofcurry.com', 'journeymart.com', 'books.google.com', 'books.google.com', 'www.whiskaffair.com', 'books.google.com', 'cities.expressindia.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'joosfood.com', 'books.google.com', 'books.google.com', 'www.hindustantimes.com', 'indfy.com', 'asiarooms.com', 'lulu.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.archanaskitchen.com', 'books.google.com', 'books.google.com', 'www.hindu.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'hebbarskitchen.com', 'www.archanaskitchen.com', 'storyofindia.com', 'www.mygingergarlickitchen.com', 'www.historyireland.com', 'books.google.com', 'www.mapsofindia.com', 'storyofindia.com', 'books.google.com', 'pepkitchen.com', 'mapsofindia.com', 'india9.com', 'articles.economictimes.indiatimes.com', 'www.silvassa-tourism.com', 'books.google.com', 'www.archanaskitchen.com', 'books.google.com', 'books.google.com', 'articles.timesofindia.indiatimes.com', 'www.indianhealthyrecipes.com', 'www.archanaskitchen.com', 'books.google.com', 'www.hindu.com', 'www.archanaskitchen.com', 'kochipost.com', 'www.archanaskitchen.com', 'indianfoodforever.com', 'mysingaporekitchen.com', 'www.whiskaffair.com', 'thediplomat.com', 'www.roymorgan.com', 'books.google.com', 'www.travellersworldwide.com', 'books.google.com', 'www.dnaindia.com', 'books.google.com', 'richindianculture.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'm.recipes.timesofindia.com', 'books.google.com', 'varadaskitchen.blogspot.com', 'www.deccanherald.com', 'sacred-texts.com', 'www.fnbnews.com', 'recipes.timesofindia.com', 'traveller.outlookindia.com', 'www.leh-ladakh-taxi-booking.com', 'www.archanaskitchen.com', 'www.deccanchronicle.com', 'books.google.com', 'books.google.com', 'www.greatbritishchefs.com', 'books.google.com', 'sacred-texts.com', 'books.google.com', 'sacred-texts.com', 'www.archanaskitchen.com', 'khanapakana.com', 'amazingarunachal.com', 'india9.com', 'articles.timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'www.indiasite.com', 'sacred-texts.com', 'thespicemess.com', 'books.google.com', 'books.google.com', 'sukhis.com', 'www.washingtonpost.com', 'books.google.com', 'food.ndtv.com', 'books.google.com', 'books.google.com', 'm.timesofindia.com', 'hindustandainik.com', 'hebbarskitchen.com', 'books.google.com', 'www.northindiancooking.com', 'sacred-texts.com', 'www.onmanorama.com', 'www.archanaskitchen.com', 'www.india-seminar.com', 'www.vegvoyages.com', 'books.google.com', 'www.streetdirectory.com', 'books.google.com', 'www.jcookingodyssey.com', 'www.blissofcooking.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'www.bhagavad-gita.org', 'asiafood.org', 'www.incredibleindia.org', 'www.bhagavad-gita.org', 'www.sahapedia.org', 'sahapedia.org', ['clinical nutrition experimental ']]",227809,Allow all users (no expiry set),163908,16 May 2003,Kaysov ,6684,6,2003-05-16,2003-05,2003
28,28,Italian-American cuisine,https://en.wikipedia.org/wiki/Italian-American_cuisine,27,0,[],[],1,0,0,18,0,0,8,0.037037037037037035,0.0,0.6666666666666666,0.0,0.0,0.037037037037037035,0,"['old.post-gazette.com', 'www.arafanelliwinery.com', 'www.delicato.com', 'www.viansa.com', 'www.winemag.com', 'scordo.com', 'foodnetwork.com', 'www.theatlantic.com', 'www.dallavallevineyards.com', 'www.rochioliwinery.com', 'www.ferrari-carano.com', 'www.aspenbusinessjournal.com', 'www.pepi.com', 'www.frankyinnewyork.com', 'www.eataly.com', 'fireflycompany.com', 'www.signorelloestate.com', 'www.pedroncelli.com', 'publishing.cdlib.org']",3644621,Allow all users (no expiry set),27268,7 January 2006,Haikupoet ,729,1,2006-01-07,2006-01,2006
29,29,British cuisine,https://en.wikipedia.org/wiki/British_cuisine,37,0,[],[],2,0,0,5,0,1,29,0.05405405405405406,0.0,0.13513513513513514,0.0,0.0,0.05405405405405406,0,"['discovernorthernireland.com', 'books.google.com', 'www.pressreader.com', 'www.india-seminar.com', 'englishbreakfastsociety.com', 'bakersfederation.org', 'www.bermuda-online.org']",7896915,Allow all users (no expiry set),19883,12 November 2006,JBull12 ,942,10,2006-11-12,2006-11,2006
30,30,Apulian cuisine,https://en.wikipedia.org/wiki/Apulian_cuisine,14,0,[],[],0,0,0,2,0,1,11,0.0,0.0,0.14285714285714285,0.0,0.0,0.0,0,"['www.tastecooking.com', 'www.gaypugliapodcast.com']",60428487,Allow all users (no expiry set),23998,6 April 2019,AlexanderVanLoon ,41,10,2019-04-06,2019-04,2019
31,31,Cuisine of Sardinia,https://en.wikipedia.org/wiki/Cuisine_of_Sardinia,2,0,[],[],1,0,0,1,0,0,0,0.5,0.0,0.5,0.0,0.0,0.5,0,"['myadventuresacrosstheworld.com', 'www.europenowjournal.org']",23475087,Allow all users (no expiry set),17909,3 July 2009,Badagnani ,40,0,2009-07-03,2009-07,2009
32,32,Lombard cuisine,https://en.wikipedia.org/wiki/Lombard_cuisine,54,0,[],[],0,0,0,1,0,0,53,0.0,0.0,0.018518518518518517,0.0,0.0,0.0,0,['www.ricetteonline.com'],32465016,Allow all users (no expiry set),44146,19 July 2011,Altes2009 ,119,1,2011-07-19,2011-07,2011
33,33,Andalusian cuisine,https://en.wikipedia.org/wiki/Andalusian_cuisine,4,0,[],[],0,0,0,2,0,0,2,0.0,0.0,0.5,0.0,0.0,0.0,0,"['www.walkingpalates.com', 'books.google.com']",3777892,Allow all users (no expiry set),5817,20 January 2006,MrDarcy ,180,2,2006-01-20,2006-01,2006
34,34,List of Jewish cuisine dishes,https://en.wikipedia.org/wiki/List_of_Jewish_cuisine_dishes,3,0,[],[],0,0,0,3,0,0,0,0.0,0.0,1.0,0.0,0.0,0.0,0,"['books.google.com', 'www.haaretz.com', 'books.google.com']",13728163,Allow all users (no expiry set),19234,14 October 2007,Tanner-Christopher ,312,0,2007-10-14,2007-10,2007
35,35,Cuisine of Liguria,https://en.wikipedia.org/wiki/Cuisine_of_Liguria,70,0,[],[],0,0,0,13,0,0,57,0.0,0.0,0.18571428571428572,0.0,0.0,0.0,0,"['www.ligucibario.com', 'www.terredilunigiana.com', 'www.ricette-tipiche.com', 'santolceseinforma.wordpress.com', 'www.ricette-tipiche.com', 'ricette.donnamoderna.com', 'www.ricette-tipiche.com', 'www.ricette-tipiche.com', 'www.ricettepercucinare.com', 'www.facebook.com', 'www.ricette-tipiche.com', 'ricette.donnamoderna.com', 'www.prodottitipici.com']",67752290,Allow all users (no expiry set),29063,24 May 2021,Spaicol ,13,2,2021-05-24,2021-05,2021
36,36,Mexican cuisine,https://en.wikipedia.org/wiki/Mexican_cuisine,107,4,"['org/10.5744/florida/9781683401674.003.0001', '10.2307/3205269', '10.1086/ahr.111.3.660', '10.3934/dcds.2015.35.1521', None, None, None, None, None, None, None, None]","[['university press of florida '], ['educational theatre journal'], ['the american historical review '], ['discrete ']]",5,0,0,28,0,1,69,0.04672897196261682,0.0,0.2616822429906542,0.037383177570093455,0.0,0.08411214953271028,4,"['www.midcitybeat.com', 'www.mexconnect.com', 'www.mexconnect.com', 'www.rickbayless.com', 'www.lasculturas.com', 'www.foxnews.com', 'www.mexconnect.com', 'www.mexconnect.com', 'www.epicurious.com', 'www.nytimes.com', 'www.mexconnect.com', 'online.wsj.com', 'www.mexconnect.com', 'www.mexconnect.com', 'www.jewishencyclopedia.com', 'www.mexiconewsnetwork.com', 'www.seriouseats.com', 'www.google.com', 'www.thedaily.com', 'gringationcancun.com', 'www.tripsavvy.com', 'issuu.com', 'mayan-yucatan-traveler.com', 'www.mexconnect.com', 'www.diariodexalapa.com', 'www.mexconnect.com', 'www.parade.com', 'www.mexconnect.com', 'ich.unesco.org', 'www.fieldmuseum.org', 'npr.org', 'www.fieldmuseum.org', 'www.laphamsquarterly.org', ['university press of florida '], ['educational theatre journal'], ['the american historical review '], ['discrete ']]",20167,Allow all users (no expiry set),80101,3 October 2001,Dmerrill ,4446,25,2001-10-03,2001-10,2001
37,37,English cuisine,https://en.wikipedia.org/wiki/English_cuisine,121,0,[],[],4,1,0,33,0,12,71,0.03305785123966942,0.008264462809917356,0.2727272727272727,0.0,0.0,0.04132231404958678,0,"['www.food.gov', 'www.januarymagazine.com', 'www.rheged.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.vegansociety.com', 'www.east-indians.com', 'www.smithsonianmag.com', 'www.pressreader.com', 'www.foodreference.com', 'www.brooklynpaper.com', 'books.google.com', 'www.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.oxforddictionaries.com', 'www.historicfood.com', 'cheftalk.com', 'books.google.com', 'www.caterersearch.com', 'www.lovefood.com', 'www.lcblondon.com', 'anglo-indianfood.blogspot.com', 'www.britishcheese.com', 'www.medievalcuisine.com', 'www.bbcamerica.com', 'www.thecaterer.com', 'www.nytimes.com', 'oed.com', 'books.google.com', 'www.india-seminar.com', 'www.menu2menu.com', 'www.european-vegetarian.org', 'icons.org', 'www.recipespastandpresent.org', 'vegsoc.org']",77208,Allow all users (no expiry set),78231,28 August 2002,62.7.21.10 ,2856,6,2002-08-28,2002-08,2002
38,38,Iranian cuisine,https://en.wikipedia.org/wiki/Iranian_cuisine,96,0,[],[],10,0,0,62,0,3,22,0.10416666666666667,0.0,0.6458333333333334,0.0,0.0,0.10416666666666667,0,"['www.reuters.com', 'books.google.com', 'ricksteves.com', 'books.google.com', 'books.google.com', 'cultureofiran.com', 'books.google.com', 'books.google.com', 'www.sfchronicle.com', 'www.huffingtonpost.com', 'books.google.com', 'books.google.com', 'www.irishtimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.cultureofiran.com', 'www.theglobeandmail.com', 'books.google.com', 'bbc.com', 'books.google.com', 'www.mehrnews.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'aashpazi.com', 'books.google.com', 'books.google.com', 'talesofakitchen.com', 'iran-daily.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'parisaskitchen.com', 'www.iranica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'bestirantravel.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'thenibble.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'electricpulp.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.iranicaonline.org', 'ostani.hamshahrilinks.org', 'faostat3.fao.org', 'www.iranicaonline.org', 'www.iran-heritage.org', 'www.iranicaonline.org', 'www.iranicaonline.org', 'www.iranicaonline.org', 'faostat.fao.org', 'www.iranicaonline.org']",2120585,Allow all users (no expiry set),62420,26 June 2005,SouthernComfort ,1875,5,2005-06-26,2005-06,2005
39,39,Egyptian cuisine,https://en.wikipedia.org/wiki/Egyptian_cuisine,43,0,[],[],5,0,0,32,0,0,6,0.11627906976744186,0.0,0.7441860465116279,0.0,0.0,0.11627906976744186,0,"['books.google.com', 'books.google.com', 'www.britannica.com', 'www.lonelyplanet.com', 'books.google.com', 'www.jonjensen.com', 'egyptian-cuisine-recipes.com', 'www.google.com', 'ribbonstopastas.com', 'books.google.com', 'www.aramcoworld.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'allrecipes.com', 'doctorfithealth.com', 'egyptbesttrip.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'allrecipes.com', 'www.bkwine.com', 'www.citylab.com', 'books.google.com', 'munchies.vice.com', 'www.atlasobscura.com', 'travelfoodatlas.com', 'books.google.com', 'www.aramcoworld.com', 'books.google.com', 'www.sbs.com', 'kew.org', 'arablit.org', 'faostat3.fao.org', 'www.reshafim.org', 'www.npr.org']",8559295,Allow all users (no expiry set),42760,22 December 2006,FunnyYetTasty ,1271,3,2006-12-22,2006-12,2006
40,40,Cuisine of Basilicata,https://en.wikipedia.org/wiki/Cuisine_of_Basilicata,86,0,[],[],0,0,0,21,0,0,65,0.0,0.0,0.2441860465116279,0.0,0.0,0.0,0,"['saporilucani.com', 'saporilucani.com', 'ricettegourmet.com', 'saporilucani.com', 'isassidimatera.com', 'www.com', 'italianroyalfood.com', 'saporilucani.com', 'fondazioneslowfood.com', 'saporilucani.com', 'saporilucani.com', 'ilsole24ore.com', 'isassidimatera.com', 'ondalucana.com', 'italianroyalfood.com', 'saporilucani.com', 'saporilucani.com', 'yumpu.com', 'foodandsoon.com', 'www.e-borghi.com', 'saporilucani.com']",69116943,Allow all users (no expiry set),40281,25 October 2021,Spaicol ,18,0,2021-10-25,2021-10,2021
41,41,Cuisine of the Indian subcontinent,https://en.wikipedia.org/wiki/Cuisine_of_the_Indian_subcontinent,4,0,[],[],0,0,0,1,0,0,3,0.0,0.0,0.25,0.0,0.0,0.0,0,['vice.com'],2687330,Allow all users (no expiry set),16453,16 September 2005,Sortan ,234,3,2005-09-16,2005-09,2005
42,42,Irish cuisine,https://en.wikipedia.org/wiki/Irish_cuisine,194,4,"['10.4000/mimmoc.1733', '10.1007/s00334-013-0417-z', '10.3318/priac.2015.115.09', None, None, None, None, None, None]","[['mémoire'], ['vegetation history and archaeobotany'], ['proceedings of the royal irish academy']]",6,1,0,13,0,0,170,0.030927835051546393,0.005154639175257732,0.06701030927835051,0.020618556701030927,0.0,0.05670103092783505,3,"['naldc.nal.usda.gov', 'www.msnbc.msn.com', 'food.com', 'www.saveur.com', 'culinarylore.com', 'www.irishtimes.com', 'www.irishtimes.com', 'galwayoysterfest.com', 'irelandseye.com', 'foodireland.com', 'www.irishtimes.com', 'www.sligoheritage.com', 'books.google.com', 'www.irishhealth.com', 'luminarium.org', 'www.worldcat.org', 'www.worldcat.org', 'journal.media-culture.org', 'www.ravensgard.org', 'www.worldcat.org', ['mémoire'], ['vegetation history and archaeobotany'], ['proceedings of the royal irish academy']]",22270189,Allow all users (no expiry set),101919,21 August 2004,Squash ,1626,1,2004-08-21,2004-08,2004
43,43,Greek cuisine,https://en.wikipedia.org/wiki/Greek_cuisine,22,1,"['10.1007/s12349-013-0123-5', None, None]",[['mediterranean journal of nutrition and metabolism']],0,0,0,2,0,0,19,0.0,0.0,0.09090909090909091,0.045454545454545456,0.0,0.045454545454545456,1,"['www.despinascafe.com', 'www.ultimate-guide-to-greek-food.com', ['mediterranean journal of nutrition and metabolism']]",12486,Allow all users (no expiry set),15670,1 November 2001,Paul Drye ,2602,12,2001-11-01,2001-11,2001
44,44,Ottoman cuisine,https://en.wikipedia.org/wiki/Ottoman_cuisine,64,2,"['10.1017/s1380203800001756', '10.1162/0022195052564252', None, None, None, None]","[['archaeological dialogues '], ['journal of interdisciplinary history ']]",0,1,0,43,0,0,18,0.0,0.015625,0.671875,0.03125,0.0,0.046875,2,"['izmir.ktb.gov', 'www.google.com', 'www.google.com', 'www.google.com', 'books.google.com', 'www.hurriyet.com', 'www.hurriyetdailynews.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.hurriyetdailynews.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.sabah.com', 'www.google.com', 'www.hurriyet.com', 'books.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.google.com', ['archaeological dialogues '], ['journal of interdisciplinary history ']]",7261681,Allow all users (no expiry set),50556,2 October 2006,OttomanReference ,301,4,2006-10-02,2006-10,2006
45,45,Neapolitan cuisine,https://en.wikipedia.org/wiki/Neapolitan_cuisine,6,0,[],[],0,0,0,1,0,0,5,0.0,0.0,0.16666666666666666,0.0,0.0,0.0,0,['foodlocate.com'],16591942,Allow all users (no expiry set),37988,26 March 2008,Guarracino ,399,0,2008-03-26,2008-03,2008
46,46,Polish cuisine,https://en.wikipedia.org/wiki/Polish_cuisine,31,0,[],[],2,0,0,8,0,0,21,0.06451612903225806,0.0,0.25806451612903225,0.0,0.0,0.06451612903225806,0,"['www.polishmeals.com', 'glosbe.com', 'books.google.com', 'www.thespruceeats.com', 'www.tastingpoland.com', 'books.google.com', 'www.beer100.com', 'www.cooksinfo.com', 'www.websters-online-dictionary.org', 'ginvodka.org']",418713,Allow all users (no expiry set),59923,3 January 2004,Halibutt ,1751,2,2004-01-03,2004-01,2004
47,47,Russian cuisine,https://en.wikipedia.org/wiki/Russian_cuisine,19,0,[],[],0,0,0,10,0,0,9,0.0,0.0,0.5263157894736842,0.0,0.0,0.0,0,"['books.google.com', 'www.advantour.com', 'enjoyyourcooking.com', 'www.pravmir.com', 'www.world-food-4u.com', 'books.google.com', 'greatbritishchefs.com', 'about.com', 'destinations.com', 'www.themoscowtimes.com']",644135,Allow all users (no expiry set),48747,9 May 2004,Marcus2 ,1425,1,2004-05-09,2004-05,2004
48,48,Albanian cuisine,https://en.wikipedia.org/wiki/Albanian_cuisine,39,1,"['10.1016/s0140-6736(97)08347-5', '9428253', None]",[['the lancet ']],6,3,0,21,0,0,10,0.15384615384615385,0.07692307692307693,0.5384615384615384,0.02564102564102564,0.0,0.2564102564102564,1,"['instat.gov', 'pdf.usaid.gov', 'usaid.gov', 'helgilibrary.com', 'www.hurriyet.com', 'books.google.com', 'scan-tv.com', 'telegrafi.com', 'www.britannica.com', 'ijoer.com', 'books.google.com', 'albaniainside.com', 'webcache.googleusercontent.com', 'telegrafi.com', 'www.britannica.com', 'drivemefoody.com', 'epicureandculture.com', 'books.google.com', 'dailysabah.com', 'books.google.com', 'webcache.googleusercontent.com', 'www.atlasobscura.com', 'books.google.com', 'books.google.com', 'agroweb.org', 'wineinstitute.org', 'anglisticum.org', 'ifama.org', 'eastagri.org', 'anglisticum.org', ['the lancet ']]",333059,Allow all users (no expiry set),38155,2 October 2003,Dori ,893,0,2003-10-02,2003-10,2003
49,49,Jewish cuisine,https://en.wikipedia.org/wiki/Jewish_cuisine,94,1,"['10.1353/jqr.0.0076', None, None]",[['the jewish quarterly review']],15,0,0,16,0,1,61,0.1595744680851064,0.0,0.1702127659574468,0.010638297872340425,0.0,0.1702127659574468,1,"['www.thespruceeats.com', 'www.thenibble.com', 'www.forward.com', 'books.google.com', 'www.haaretz.com', 'www.jewishencyclopedia.com', 'forward.com', 'net.com', 'momentmag.com', 'www.bbc.com', 'about.com', 'www.nytimes.com', 'jewishlinknj.com', 'www.elitetraveler.com', 'www.kosher.com', 'www.huffingtonpost.com', 'bckosher.org', 'www.jewishvirtuallibrary.org', 'www.crcweb.org', 'www.asor.org', 'www.chabad.org', 'www.jewishvirtuallibrary.org', 'www.mechon-mamre.org', 'www.chabad.org', 'www.chabad.org', 'www.jewishvirtuallibrary.org', 'www.mechon-mamre.org', 'www.jewishvirtuallibrary.org', 'stories.thejewishmuseum.org', 'www.chabad.org', 'www.chabad.org', ['the jewish quarterly review']]",1290526,Allow all users (no expiry set),63582,17 December 2004,Saintswithin ,1614,1,2004-12-17,2004-12,2004
50,50,Mongolian cuisine,https://en.wikipedia.org/wiki/Mongolian_cuisine,10,0,[],[],0,0,0,1,0,0,9,0.0,0.0,0.1,0.0,0.0,0.0,0,['www.behindcity.com'],5571891,Allow all users (no expiry set),12305,15 June 2006,Latebird ,464,0,2006-06-15,2006-06,2006
51,51,Du fait de cuisine,https://en.wikipedia.org/wiki/Du_fait_de_cuisine,2,0,[],[],0,0,0,0,0,0,2,0.0,0.0,0.0,0.0,0.0,0.0,0,[],24227321,Allow all users (no expiry set),817,5 September 2009,Wetman ,21,7,2009-09-05,2009-09,2009
52,52,Cypriot cuisine,https://en.wikipedia.org/wiki/Cypriot_cuisine,4,0,[],[],0,0,0,2,0,0,2,0.0,0.0,0.5,0.0,0.0,0.0,0,"['www.travelerslunchbox.com', 'www.visitcyprus.com']",2582022,Allow all users (no expiry set),21282,31 August 2005,195.14.141.58 ,658,5,2005-08-31,2005-08,2005
53,53,Italian Eritrean cuisine,https://en.wikipedia.org/wiki/Italian_Eritrean_cuisine,4,0,[],[],0,0,0,3,0,0,1,0.0,0.0,0.75,0.0,0.0,0.0,0,"['books.google.com', 'www.washingtoncitypaper.com', 'asmarabrewery.com']",32125586,Allow all users (no expiry set),4563,18 June 2011,Hidudes1000 ,47,0,2011-06-18,2011-06,2011
54,54,Icelandic cuisine,https://en.wikipedia.org/wiki/Icelandic_cuisine,6,0,[],[],0,0,0,1,0,0,5,0.0,0.0,0.16666666666666666,0.0,0.0,0.0,0,['www.newyorker.com'],5642461,Allow all users (no expiry set),35966,20 June 2006,Green caterpillar ,563,1,2006-06-20,2006-06,2006
55,55,Dutch cuisine,https://en.wikipedia.org/wiki/Dutch_cuisine,19,0,[],[],4,0,0,7,0,0,8,0.21052631578947367,0.0,0.3684210526315789,0.0,0.0,0.21052631578947367,0,"['books.google.com', 'www.thehollandring.com', 'www.web-books.com', 'thedutchtable.com', 'holland.com', 'books.google.com', 'about.com', 'aboutus.org', 'www.dbnl.org', 'www.culinaryhistoriansny.org', 'www.sca-indo.org']",918733,Allow all users (no expiry set),55859,21 August 2004,Squash ,1655,16,2004-08-21,2004-08,2004
56,56,Iraqi cuisine,https://en.wikipedia.org/wiki/Iraqi_cuisine,33,1,"['10.1016/s0262-1762(10)70355-2', None, None]",[['world pumps']],3,0,0,15,0,0,14,0.09090909090909091,0.0,0.45454545454545453,0.030303030303030304,0.0,0.12121212121212122,1,"['blog.foodpairing.com', 'www.tasteofbeirut.com', 'www.saudiaramcoworld.com', 'www.hungrypaprikas.com', 'www.kosher.com', 'www.internationalcuisine.com', 'www.smithakalluraya.com', 'books.google.com', 'www.al-monitor.com', 'www.indianhealthyrecipes.com', 'www.thingsasian.com', 'latimesblogs.latimes.com', 'books.google.com', 'justgotochef.com', 'www.bbc.com', 'www.laphamsquarterly.org', 'historyetc.org', 'etc.worldhistory.org', ['world pumps']]",2322115,Allow all users (no expiry set),35547,27 July 2005,81.153.74.21 ,1156,1,2005-07-27,2005-07,2005
57,57,Bangladeshi cuisine,https://en.wikipedia.org/wiki/Bangladeshi_cuisine,19,0,[],[],0,0,0,11,0,2,6,0.0,0.0,0.5789473684210527,0.0,0.0,0.0,0,"['www.withaspin.com', 'books.google.com', 'www.daily-sun.com', 'www.daily-sun.com', 'blogs.wsj.com', 'www.daily-sun.com', 'www.localguidesconnect.com', 'archive.dhakatribune.com', 'offroadbangladesh.com', 'www.nytimes.com', 'www.foodiez.com']",3011692,Allow all users (no expiry set),16123,27 October 2005,Aloodum ,1005,0,2005-10-27,2005-10,2005
58,58,Portuguese cuisine,https://en.wikipedia.org/wiki/Portuguese_cuisine,81,1,"['10.1080/14664650500314513', None, None]",[['american nineteenth century history ']],4,6,0,32,0,0,38,0.04938271604938271,0.07407407407407407,0.3950617283950617,0.012345679012345678,0.0,0.13580246913580246,1,"['tradicional.dgadr.gov', 'tradicional.dgadr.gov', 'tradicional.dgadr.gov', 'tradicional.dgadr.gov', 'tradicional.dgadr.gov', 'tradicional.dgadr.gov', 'www.vogue.com', 'books.google.com', 'www.bikeonelas.com', 'brill.com', 'wetravelportugal.com', 'books.google.com', 'www.google.com', 'www.amasscook.com', 'www.amasscook.com', 'www.lalanguefrancaise.com', 'thestar.com', 'bbc.com', 'www.internationalcuisine.com', 'books.google.com', 'newstatesman.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'www.portugalthings.com', 'kidbite.wordpress.com', 'www.portaldojardim.com', 'www.aaronokada.com', 'www.bol.com', 'www.topdeportugal.com', 'books.google.com', 'www.gloriascafe.com', 'filter.com', 'seattle.eater.com', 'www.smh.com', 'www.forbes.com', 'kyotofoodie.com', 'igbp-portugal.org', 'smithsonianassociates.org', 'ourworldindata.org', 'dicionario.priberam.org', ['american nineteenth century history ']]",918711,Allow all users (no expiry set),58218,21 August 2004,Squash ,1585,16,2004-08-21,2004-08,2004
59,59,Serbian cuisine,https://en.wikipedia.org/wiki/Serbian_cuisine,15,0,[],[],1,1,0,6,0,0,7,0.06666666666666667,0.06666666666666667,0.4,0.0,0.0,0.13333333333333333,0,"['www.zis.gov', 'www.lonelyplanet.com', 'www.balkanfoodrecipes.com', 'www.vreme.com', 'kuhinjica.forumotion.com', 'www.ekapija.com', 'sputnik-news.com', 'www.gmo-free-regions.org']",2015602,Allow all users (no expiry set),32770,9 June 2005,213.240.13.238 ,1155,4,2005-06-09,2005-06,2005
60,60,Udupi cuisine,https://en.wikipedia.org/wiki/Udupi_cuisine,9,0,[],[],0,0,0,6,0,0,3,0.0,0.0,0.6666666666666666,0.0,0.0,0.0,0,"['www.thehinduonnet.com', 'www.in.rediff.com', 'mumbaimirror.com', 'www.udupitourism.com', 'udupi-recipes.com', 'www.karnataka.com']",3560438,Allow all users (no expiry set),12041,29 December 2005,Balaji Varma ,443,3,2005-12-29,2005-12,2005
61,61,New American cuisine,https://en.wikipedia.org/wiki/New_American_cuisine,5,0,[],[],0,0,0,2,0,0,3,0.0,0.0,0.4,0.0,0.0,0.0,0,"['philipmarie.com', 'www.abebooks.com']",4604855,Allow all users (no expiry set),2408,2 April 2006,Haikupoet ,72,0,2006-04-02,2006-04,2006
62,62,Norwegian cuisine,https://en.wikipedia.org/wiki/Norwegian_cuisine,9,0,[],[],1,0,0,3,0,0,5,0.1111111111111111,0.0,0.3333333333333333,0.0,0.0,0.1111111111111111,0,"['www.norwegianamerican.com', 'www.bbc.com', 'www.visitnorway.com', 'www.worldcat.org']",2215144,Allow all users (no expiry set),29096,11 July 2005,Vikingstad ,866,3,2005-07-11,2005-07,2005
63,63,American Chinese cuisine,https://en.wikipedia.org/wiki/American_Chinese_cuisine,71,2,"['10.1016/j.ijhm.2008.10.008', '10.1093/acrefore/9780199329175.013.273', None, None, None, None]","[['international journal of hospitality management '], ['oxford research encyclopedia ']]",8,1,0,45,0,0,15,0.11267605633802817,0.014084507042253521,0.6338028169014085,0.028169014084507043,0.0,0.15492957746478872,2,"['factfinder.census.gov', 'fromaway.com', 'www.philly.com', 'www.thehindu.com', 'www.smithsonianmag.com', 'www.nytimes.com', 'www.nyfoodstory.com', 'cnneatocracy.wordpress.com', 'about.com', 'www.nytimes.com', 'www.nytimes.com', 'radiichina.com', 'www.vice.com', 'www.wsj.com', 'chow.com', 'huffingtonpost.com', 'news.asianweek.com', 'books.google.com', 'www.nytimes.com', 'www.thespruceeats.com', 'www.ming.com', 'www.theodysseyonline.com', 'www.latimes.com', 'thaitable.com', 'www.latimes.com', 'theatlantic.com', 'luckypeach.com', 'queensbuzz.com', 'about.com', 'www.nytimes.com', 'canyoustayfordinner.com', 'radiichina.com', 'www.nytimes.com', 'www.nytimes.com', 'books.google.com', 'www.latimes.com', 'www.haaretz.com', 'www.scoutingny.com', 'rasamalaysia.com', 'www.nytimes.com', 'www.pandarg.com', 'www.nytimes.com', 'www.insider.com', 'food.com', 'www.nytimes.com', 'imdiversity.com', 'asian-studies.org', 'www.pri.org', 'www.npr.org', 'www.jstor.org', 'www.scpr.org', 'www.npr.org', 'www.newuniversity.org', 'cambridgehistory.org', ['international journal of hospitality management '], ['oxford research encyclopedia ']]",1558,Allow all users (no expiry set),53914,5 November 2001,24.4.254.xxx ,1813,0,2001-11-05,2001-11,2001
64,64,Pie in American cuisine,https://en.wikipedia.org/wiki/Pie_in_American_cuisine,73,0,[],[],4,3,0,65,0,0,1,0.0547945205479452,0.0410958904109589,0.8904109589041096,0.0,0.0,0.0958904109589041,0,"['blogs.loc.gov', 'www.maine.gov', 'history.nebraska.gov', 'www.newspapers.com', 'www.newspapers.com', 'www.newspapers.com', 'www.google.com', 'www.newspapers.com', 'www.newspapers.com', 'cooking.nytimes.com', 'www.newspapers.com', 'www.newspapers.com', 'www.newspapers.com', 'www.google.com', 'www.newspapers.com', 'www.southernliving.com', 'www.newspapers.com', 'www.google.com', 'www.newspapers.com', 'www.newspapers.com', 'www.newspapers.com', 'www.google.com', 'www.newspapers.com', 'www.latimes.com', 'www.nhmagazine.com', 'www.newspapers.com', 'www.youtube.com', 'www.newspapers.com', 'www.newspapers.com', 'www.heraldnews.com', 'www.newspapers.com', 'www.newspapers.com', 'www.newspapers.com', 'www.newspapers.com', 'www.southernliving.com', 'www.newspapers.com', 'www.google.com', 'www.newspapers.com', 'www.newspapers.com', 'www.chicagotribune.com', 'www.newspapers.com', 'www.newspapers.com', 'www.newspapers.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.newspapers.com', 'www.newspapers.com', 'www.newspapers.com', 'www.newspapers.com', 'www.newspapers.com', 'www.newspapers.com', 'www.newspapers.com', 'www.newenglandhistoricalsociety.com', 'www.tasteofhome.com', 'www.newspapers.com', 'www.newspapers.com', 'www.newspapers.com', 'www.southernliving.com', 'www.newspapers.com', 'www.newspapers.com', 'www.google.com', 'www.newspapers.com', 'www.google.com', 'www.newspapers.com', 'www.google.com', 'www.newspapers.com', 'www.southernliving.com', 'www.piecouncil.org', 'www.piecouncil.org', 'alfafarmers.org', 'dictionary.cambridge.org']",65542369,Allow all users (no expiry set),41465,9 October 2020,Spudlace ,112,1,2020-10-09,2020-10,2020
65,65,Kurdish cuisine,https://en.wikipedia.org/wiki/Kurdish_cuisine,11,0,[],[],3,0,0,7,0,1,0,0.2727272727272727,0.0,0.6363636363636364,0.0,0.0,0.2727272727272727,0,"['www.youtube.com', 'cuisinemiddleast.com', 'www.youtube.com', 'cuisinemiddleast.com', 'cache:eq_abt_wv48j:www.saradistribution.com', 'bestofvegan.com', 'kurdishbike.com', 'krg.org', 'krg.org', 'bnk.institutkurde.org']",3912255,Allow all users (no expiry set),12826,31 January 2006,Diyako ,256,0,2006-01-31,2006-01,2006
66,66,Armenian cuisine,https://en.wikipedia.org/wiki/Armenian_cuisine,72,6,"['10.1016/b978-0-12-394801-4.00026-0', '10.1016/j.jef.2016.05.005', '10.1016/b978-0-444-63666-9.00008-x', '10.1016/j.jef.2016.01.003', '10.1016/j.smallrumres.2011.09.021', '10.1016/b978-0-12-800850-8.00001-6', None, None, None, None, None, None, None, None, None, None, None, None]","[[' elsevier'], [' journal of ethnic foods'], [' elsevier'], [' journal of ethnic foods'], [' small ruminant research'], [' academic press']]",6,0,0,30,0,1,29,0.08333333333333333,0.0,0.4166666666666667,0.08333333333333333,0.0,0.16666666666666666,6,"['books.google.com', 'www.road-to-armenia.com', 'www.topliquor.com', 'www.armenianow.com', 'www.milliyet.com', 'heghineh.com', 'books.google.com', 'articles.latimes.com', 'books.google.com', 'books.google.com', 'answers.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.smithsonianmag.com', 'www.sozcu.com', 'www.kanald.com', 'www.bostonglobe.com', 'books.google.com', 'books.google.com', 'cooking.nytimes.com', 'www.youtube.com', 'www.oxfordreference.com', 'www.tacentral.com', 'www.travelchannel.com', 'www.jdemirdjian.com', 'www.sptimes.com', 'www.chowhound.com', 'www.houshamadyan.org', 'www.houshamadyan.org', 'www.houshamadyan.org', 'www.houshamadyan.org', 'fita.org', 'www.saintsarkis.org', [' elsevier'], [' journal of ethnic foods'], [' elsevier'], [' journal of ethnic foods'], [' small ruminant research'], [' academic press']]",6582433,Allow all users (no expiry set),66338,20 August 2006,Eupator ,1018,12,2006-08-20,2006-08,2006
67,67,History of Indian cuisine,https://en.wikipedia.org/wiki/History_of_Indian_cuisine,77,7,"['10.1371/journal.pone.0073682', '10.1038/srep19157', '10.1086/383236', '10.1086/658860', '10.1086/318200', '10.1371/journal.pone.0095714', '10.1017/s0003598x00048249', '24040024', '26754573', '15077202', None, '11133362', '24806472', None, '3770703', '4709632', '1181978', None, '1235289', '4012948', None]","[['plos one '], ['scientific reports '], [' am j hum genet '], [' curr anthropol '], [' am j hum genet '], ['plos one '], [' antiquity ']]",3,2,0,42,0,0,24,0.03896103896103896,0.025974025974025976,0.5454545454545454,0.09090909090909091,0.0,0.15584415584415584,7,"['food.gov', 'www.food.gov', 'books.google.com', 'books.google.com', 'asiarooms.com', 'hindustandainik.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.bestindianfoodcatering.com', 'www.livemint.com', 'books.google.com', 'books.google.com', 'rediff.com', 'www.asianage.com', 'books.google.com', 'www.globalpost.com', 'books.google.com', 'timesofindia.indiatimes.com', 'brill.com', 'server2.docfoc.com', 'www.history.com', 'books.google.com', 'www.washingtonpost.com', 'theculturetrip.com', 'timesofindia.indiatimes.com', 'www.travellersworldwide.com', 'slate.com', 'www.hindustantimes.com', 'about.com', 'economictimes.indiatimes.com', 'brill.com', 'www.vegvoyages.com', 'archaeology.about.com', 'books.google.com', 'www.esamskriti.com', 'www.washingtonpost.com', 'vice.com', 'books.google.com', 'www.india-seminar.com', 'books.google.com', 'www.streetdirectory.com', 'www.nytimes.com', 'www.pri.org', 'www.pri.org', 'whc.unesco.org', ['plos one '], ['scientific reports '], [' am j hum genet '], [' curr anthropol '], [' am j hum genet '], ['plos one '], [' antiquity ']]",17837671,Allow all users (no expiry set),41007,8 June 2008,Shyamsunder ,144,1,2008-06-08,2008-06,2008
68,68,Welsh cuisine,https://en.wikipedia.org/wiki/Welsh_cuisine,54,0,[],[],0,2,0,36,0,0,16,0.0,0.037037037037037035,0.6666666666666666,0.0,0.0,0.037037037037037035,0,"['food.gov', 'www.food.gov', 'infoweb.newsbank.com', 'tynant.com', 'literati.credoreference.com', 'books.google.com', 'books.google.com', 'books.google.com', 'infoweb.newsbank.com', 'www.sparknotes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'literati.credoreference.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'literati.credoreference.com', 'books.google.com', 'literati.credoreference.com', 'books.google.com', 'princesgate.com', 'literati.credoreference.com', 'books.google.com', 'literati.credoreference.com', 'books.google.com']",50034045,Allow all users (no expiry set),43375,7 July 2005,Wikisurfer1 ,645,0,2005-07-07,2005-07,2005
69,69,Assamese cuisine,https://en.wikipedia.org/wiki/Assamese_cuisine,10,1,"['10.1016/j.dit.2013.09.002', None, None]",[['drug invention today ']],0,0,0,4,0,0,5,0.0,0.0,0.4,0.1,0.0,0.1,1,"['www.india-seminar.com', 'www.uppercrustindia.com', 'recipes.timesofindia.com', 'time.com', ['drug invention today ']]",1810291,Allow all users (no expiry set),24847,28 April 2005,Chaipau ,833,2,2005-04-28,2005-04,2005
70,70,Lithuanian cuisine,https://en.wikipedia.org/wiki/Lithuanian_cuisine,38,1,[],[],1,0,0,6,0,0,30,0.02631578947368421,0.0,0.15789473684210525,0.02631578947368421,0.0,0.05263157894736842,0,"['www.food.com', 'kulinarinispaveldas.blogspot.com', 'kulinarinispaveldas.blogspot.com', 'curioustovisit.com', 'www.thelatinlibrary.com', 'youtube.com', 'www.brewersofeurope.org']",948976,Allow all users (no expiry set),64452,1 September 2004,Kpjas ,934,1,2004-09-01,2004-09,2004
71,71,Vegetarian cuisine,https://en.wikipedia.org/wiki/Vegetarian_cuisine,10,3,"['10.1017/s000711451400261x', '10.1079/pns2005481', '10.2337/dc10-1221', None, '16441942', '21411506', '4232985', None, '3114510']","[['british journal of nutrition'], ['proceedings of the nutrition society'], ['diabetes care']]",3,1,0,1,0,0,2,0.3,0.1,0.1,0.3,0.0,0.7,3,"['www.nhlbi.nih.gov', 'www.healthline.com', 'www.mayoclinic.org', 'www.vegsoc.org', 'ivu.org', ['british journal of nutrition'], ['proceedings of the nutrition society'], ['diabetes care']]",32601,Allow all users (no expiry set),24188,29 September 2001,65.31.133.xxx ,748,2,2001-09-29,2001-09,2001
72,72,Scottish cuisine,https://en.wikipedia.org/wiki/Scottish_cuisine,19,0,[],[],0,0,0,6,0,0,13,0.0,0.0,0.3157894736842105,0.0,0.0,0.0,0,"['news.google.com', 'www.edinburghnews.scotsman.com', 'www.historichighlanders.com', 'www.geraldeneholt.com', 'www.radiotimes.com', 'www.taste-of-scotland.com']",6169255,Allow all users (no expiry set),21698,29 July 2006,Nach0king ,1100,2,2006-07-29,2006-07,2006
73,73,Israeli cuisine,https://en.wikipedia.org/wiki/Israeli_cuisine,134,1,"['10.1177/1468796813519428', None, None]",[[' ethnicities']],6,0,0,31,0,0,96,0.04477611940298507,0.0,0.23134328358208955,0.007462686567164179,0.0,0.05223880597014925,1,"['library-genesis.com', 'www.myjewishlearning.com', 'books.google.com', 'ynetnews.com', 'thejc.com', 'www.the-eucalyptus.com', 'dancingcamel.com', 'www.gemsinisrael.com', 'www.themarker.com', 'ynetnews.com', 'www.jpost.com', 'www.ynetnews.com', 'blogs.forward.com', 'www.ynetnews.com', 'www.winebusiness.com', 'www.myjewishlearning.com', 'www.haaretz.com', 'www.foxnews.com', 'www.virtualjerusalem.com', 'www.haaretz.com', 'www.haaretz.com', 'books.google.com', 'halachipedia.com', 'www.strauss-group.com', 'www.myjewishlearning.com', 'www.nytimes.com', 'www.haaretz.com', 'forward.com', 'www.encyclopedia.com', 'www.israel-travel-tips.com', 'www.myjewishlearning.com', 'www.israel21c.org', 'www.israel21c.org', 'www.jewishvirtuallibrary.org', 'www.jewishvirtuallibrary.org', 'www.jewishvirtuallibrary.org', 'faostat3.fao.org', [' ethnicities']]",11447140,Require extended confirmed access (no expiry set),88965,27 May 2007,Acidburn24m ,1721,1,2007-05-27,2007-05,2007
74,74,Romanian cuisine,https://en.wikipedia.org/wiki/Romanian_cuisine,27,0,[],[],2,0,0,12,0,0,13,0.07407407407407407,0.0,0.4444444444444444,0.0,0.0,0.07407407407407407,0,"['www.cooks.com', 'www.exploringromania.com', 'www.huffingtonpost.com', 'www.vulpeabucatar.com', 'filter.com', 'www.roconsulboston.com', 'www.pbase.com', 'www.kitchencookingrecipes.com', 'educations.com', 'www.imperialtransilvania.com', 'www.regard-est.com', 'family.webshots.com', 'www.ivu.org', 'faostat.fao.org']",1245931,Allow all users (no expiry set),32343,5 December 2004,Bogdangiusca ,1052,3,2004-12-05,2004-12,2004
75,75,History of Chinese cuisine,https://en.wikipedia.org/wiki/History_of_Chinese_cuisine,80,0,[],[],1,0,0,19,0,0,60,0.0125,0.0,0.2375,0.0,0.0,0.0125,0,"['books.google.com', 'books.google.com', 'books.google.com', 'www.chinapage.com', 'books.google.com', 'books.google.com', 'books.google.com', 'food52.com', 'books.google.com', 'books.google.com', 'www.yhnkzq.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.worldcat.org']",3949800,Allow all users (no expiry set),50079,3 February 2006,Ram32110 ,619,2,2006-02-03,2006-02,2006
76,76,Pakistani cuisine,https://en.wikipedia.org/wiki/Pakistani_cuisine,25,0,[],[],1,0,0,15,0,0,9,0.04,0.0,0.6,0.0,0.0,0.04,0,"['dominos.com', 'pakistantumhetoho.com', 'www.thehindu.com', 'sindhikhazana.com', 'nation.com', 'www.pizzahut.com', 'www.papajohns.com', 'www.curryflow.com', 'www.papajohns.com', 'www.kfcpakistan.com', 'bawarchi.com', 'mcdonalds.com', 'www.subway.com', 'www.sairamtour.com', 'www.dunkindonuts.com', 'jn.nutrition.org']",429283,Allow all users (no expiry set),37126,13 January 2004,DigiBullet ,2076,6,2004-01-13,2004-01,2004
77,77,Ancient Roman cuisine,https://en.wikipedia.org/wiki/Ancient_Roman_cuisine,52,2,"['10.1017/cbo9780511585395', '10.2752/155280105778055407', None, None, None, None]","[['cambridge university press'], ['food']]",0,0,0,4,0,0,46,0.0,0.0,0.07692307692307693,0.038461538461538464,0.0,0.038461538461538464,2,"['books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', ['cambridge university press'], ['food']]",214980,Allow all users (no expiry set),30588,23 April 2003,Junesun ,2134,5,2003-04-23,2003-04,2003
78,78,St. Louis cuisine,https://en.wikipedia.org/wiki/St._Louis_cuisine,8,0,[],[],0,0,0,4,0,0,4,0.0,0.0,0.5,0.0,0.0,0.0,0,"['ksdk.com', 'explorestlouis.com', 'www.mamasonthehill.com', 'books.google.com']",41569450,Allow all users (no expiry set),6027,7 January 2014,Kazvorpal ,267,0,2014-01-07,2014-01,2014
79,79,Outline of cuisines,https://en.wikipedia.org/wiki/Outline_of_cuisines,9,0,[],[],1,0,0,5,0,1,2,0.1111111111111111,0.0,0.5555555555555556,0.0,0.0,0.1111111111111111,0,"['www.britannica.com', 'hadithcollection.com', 'www.ldoceonline.com', 'hadithcollection.com', 'books.google.com', 'dictionary.cambridge.org']",39466243,Allow all users (no expiry set),12731,23 May 2013,The Transhumanist ,84,0,2013-05-23,2013-05,2013
80,80,Modernist Cuisine,https://en.wikipedia.org/wiki/Modernist_Cuisine,25,0,[],[],3,0,0,21,0,0,1,0.12,0.0,0.84,0.0,0.0,0.12,0,"['www.bloomberg.com', 'eater.com', 'www.forbes.com', 'www.bloomberg.com', 'www.latimes.com', 'old.cookbookfair.com', 'modernistcuisine.com', 'www.cookbookfair.com', 'www.nytimes.com', 'www.google.com', 'www.popsci.com', 'modernistcuisine.com', 'www.featureshoot.com', 'intellectualventures.com', 'www.wired.com', 'modernistcuisine.com', 'amazon.com', 'www.saveur.com', 'modernistcuisine.com', 'www.wsj.com', 'www.newyorker.com', 'www.pacificsciencecenter.org', 'www.jamesbeard.org', 'www.worldcat.org']",31637084,Allow all users (no expiry set),17752,30 April 2011,Stefan-S ,158,2,2011-04-30,2011-04,2011
81,81,Bosnia and Herzegovina cuisine,https://en.wikipedia.org/wiki/Bosnia_and_Herzegovina_cuisine,4,0,[],[],0,0,0,1,0,0,3,0.0,0.0,0.25,0.0,0.0,0.0,0,['sbs.com'],5668862,Allow all users (no expiry set),10189,22 June 2006,DJ Bungi ,800,1,2006-06-22,2006-06,2006
82,82,Circassian cuisine,https://en.wikipedia.org/wiki/Circassian_cuisine,4,0,[],[],0,0,0,4,0,0,0,0.0,0.0,1.0,0.0,0.0,0.0,0,"['www.youtube.com', 'www.circassianworld.com', 'www.circassianworld.com', 'www.youtube.com']",39935792,Allow all users (no expiry set),10315,11 July 2013,Samizambak ,111,0,2013-07-11,2013-07,2013
83,83,Jharkhandi cuisine,https://en.wikipedia.org/wiki/Jharkhandi_cuisine,18,0,[],[],1,0,0,16,0,0,1,0.05555555555555555,0.0,0.8888888888888888,0.0,0.0,0.05555555555555555,0,"['pandareviewz.com', 'www.telegraphindia.com', 'indianvagabond.com', 'www.telegraphindia.com', 'www.telegraphindia.com', 'zeenews.india.com', 'books.google.com', 'www.telegraphindia.com', 'economictimes.indiatimes.com', 'books.google.com', 'www.thehindu.com', 'www.telegraphindia.com', 'www.inuth.com', 'books.google.com', 'cookpad.com', 'www.bhoomika.com', 'www.jharkhandtourism.org']",15689741,Allow all users (no expiry set),10265,10 February 2008,Kachhapbk2 ,285,6,2008-02-10,2008-02,2008
84,84,Sylheti cuisine,https://en.wikipedia.org/wiki/Sylheti_cuisine,46,0,[],[],2,0,0,32,0,2,10,0.043478260869565216,0.0,0.6956521739130435,0.0,0.0,0.043478260869565216,0,"['www.prothomalo.com', 'archive.prothom-alo.com', 'www.aljazeera.com', 'www.bd-journal.com', 'www.thestatesman.com', 'www.ntvbd.com', 'www.breadexperience.com', 'archive1.ittefaq.com', 'indianexpress.com', 'www.historic-uk.com', 'www.sylheterdak.com', 'bangladeshiweus.com', 'sylheterdak.com', 'www.jugantor.com', 'www.mid-day.com', 'www.ft.com', 'web.dailyjanakantha.com', 'www.sciencedaily.com', 'www.bhorerkagoj.com', 'frontline.thehindu.com', 'jalalabadbarta.com', 'www.daily-sun.com', 'thehindubusinessline.com', 'www.banglatribune.com', 'books.google.com', 'banglanews24.com', 'bdnews24.com', 'www.greatbritishchefs.com', 'www.prothomalo.com', 'khadizaskitchen.com', 'www.atlasobscura.com', 'www.uniindia.com', 'npr.org', 'www.sahapedia.org']",63766442,Allow all users (no expiry set),25020,25 April 2020,AbuSayeed ,55,0,2020-04-25,2020-04,2020
85,85,Cuisine of Dorset,https://en.wikipedia.org/wiki/Cuisine_of_Dorset,15,0,[],[],0,0,0,0,0,0,15,0.0,0.0,0.0,0.0,0.0,0.0,0,[],24561462,Allow all users (no expiry set),7849,3 October 2009,MasterOfHisOwnDomain ,62,1,2009-10-03,2009-10,2009
86,86,Note by Note cuisine,https://en.wikipedia.org/wiki/Note_by_Note_cuisine,5,1,"['10.1186/2044-7248-2-1', None, None]",[['flavour ']],1,0,0,0,0,0,3,0.2,0.0,0.0,0.2,0.0,0.4,1,"['www.pbs.org', ['flavour ']]",41031835,Allow all users (no expiry set),11879,9 November 2013,Tentinator ,26,0,2013-11-09,2013-11,2013
87,87,Cuisine of Ceredigion,https://en.wikipedia.org/wiki/Cuisine_of_Ceredigion,85,0,[],[],1,0,0,3,0,0,81,0.011764705882352941,0.0,0.03529411764705882,0.0,0.0,0.011764705882352941,0,"['www.gunsonpegs.com', 'www.finewaters.com', 'www.gunsonpegs.com', 'www.nationaltrust.org']",56164461,Allow all users (no expiry set),43516,29 December 2017,Vouliagmeni ,86,0,2017-12-29,2017-12,2017
88,88,Cuisine of Monmouthshire,https://en.wikipedia.org/wiki/Cuisine_of_Monmouthshire,113,0,[],[],4,0,0,8,0,0,101,0.035398230088495575,0.0,0.07079646017699115,0.0,0.0,0.035398230088495575,0,"['www.madeinmonmouthshire.com', 'www.visitmonmouthshire.com', 'britainssecrettreasures.blogspot.com', 'www.bbc.com', 'www.abergavennychronicle.com', 'www.visitmonmouthshire.com', 'www.bbc.com', 'www.cidercellars.com', 'friendsoffriendlesschurches.org', 'www.sustainweb.org', 'www.gwentwildlife.org', 'www.gwentwildlife.org']",62161487,Allow all users (no expiry set),63499,25 October 2019,Vouliagmeni ,48,0,2019-10-25,2019-10,2019
89,89,Cuisine of Pembrokeshire,https://en.wikipedia.org/wiki/Cuisine_of_Pembrokeshire,64,0,[],[],3,0,0,1,0,1,59,0.046875,0.0,0.015625,0.0,0.0,0.046875,0,"['www.visitwales.com', 'bumblebeeconservation.org', 'vegetarianforlife.org', 'www.pembrokeshire.camra.org']",51548076,Allow all users (no expiry set),37773,8 September 2016,Vouliagmeni ,85,0,2016-09-08,2016-09,2016
90,90,Pottage,https://en.wikipedia.org/wiki/Pottage,15,0,[],[],0,0,0,4,0,1,10,0.0,0.0,0.26666666666666666,0.0,0.0,0.0,0,"['books.google.com', 'books.google.com', 'www.dailytrust.com', 'books.google.com']",10955928,Allow all users (no expiry set),11935,28 April 2007,Elrith ,175,0,2007-04-28,2007-04,2007
91,91,Le Viandier,https://en.wikipedia.org/wiki/Le_Viandier,5,0,[],[],0,0,0,1,0,0,4,0.0,0.0,0.2,0.0,0.0,0.0,0,['books.google.com'],3398583,Allow all users (no expiry set),5629,12 December 2005,TomPurdue ,76,0,2005-12-12,2005-12,2005
92,92,Lancelot de Casteau,https://en.wikipedia.org/wiki/Lancelot_de_Casteau,3,0,[],[],0,0,0,2,0,0,1,0.0,0.0,0.6666666666666666,0.0,0.0,0.0,0,"['books.google.com', 'www.amazon.com']",34732474,Allow all users (no expiry set),3159,14 February 2012,Macrakis ,27,0,2012-02-14,2012-02,2012
93,93,List of desserts,https://en.wikipedia.org/wiki/List_of_desserts,4,0,[],[],0,0,0,3,0,0,1,0.0,0.0,0.75,0.0,0.0,0.0,0,"['books.google.com', 'www.britannica.com', 'www.merriam-webster.com']",41535911,Allow all users (no expiry set),46778,3 January 2014,Northamerica1000 ,725,7,2014-01-03,2014-01,2014
94,94,Food history,https://en.wikipedia.org/wiki/Food_history,43,4,"['10.1163/187247111x579296', '10.1017/s0026749x00013627', '10.1093/qje/qjr009', None, None, '22073408', None, None, None]","[['european journal of jewish studies'], ['modern asian studies'], [' [[quarterly journal of economics']]",3,1,0,4,0,0,31,0.06976744186046512,0.023255813953488372,0.09302325581395349,0.09302325581395349,0.0,0.18604651162790697,3,"['plants.usda.gov', 'books.google.com', 'books.google.com', 'books.google.com', 'www.myjewishlearning.com', 'libcom.org', 'foodtimeline.org', 'www.nypl.org', ['european journal of jewish studies'], ['modern asian studies'], [' [[quarterly journal of economics']]",21955305,Allow all users (no expiry set),36577,13 March 2009,SimonP ,420,1,2009-03-13,2009-03,2009
95,95,Squab,https://en.wikipedia.org/wiki/Squab,57,9,"['10.1186/s42779-020-00053-5', '10.1525/gfc.2005.5.2.50', '10.1525/gfc.2009.9.1.36', '10.3382/ps.2008-00217', '10.1093/ps/80.1.66', '10.1186/1297-9686-24-6-553', '10.1525/gfc.2004.4.4.25', '10.1093/oxfordjournals.jhered.a111314', '10.1901/jeab.1986.45-229', None, None, None, '19439644', '11214338', None, None, None, '3958668', None, None, None, None, None, '2711175', None, None, '1348231']","[['journal of ethnic foods'], ['[[gastronomica'], ['gastronomica'], ['poultry science '], ['poultry science'], [' genetics selection evolution '], ['gastronomica'], ['[[journal of heredity'], ['journal of the experimental analysis of behavior']]",3,1,0,21,0,2,21,0.05263157894736842,0.017543859649122806,0.3684210526315789,0.15789473684210525,0.0,0.22807017543859648,9,"['www.dpi.nsw.gov', 'books.google.com', 'books.google.com', 'books.google.com', 'arfjournals.com', 'www.nytimes.com', 'books.google.com', 'books.google.com', 'events.nytimes.com', 'www.holidify.com', 'www.greatitalianchefs.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.eastmojo.com', 'www.cnngo.com', 'www.outlookindia.com', 'www.theage.com', 'www.allqdup.com', 'www.firstpost.com', 'm.timesofindia.com', 'www.qualitativesociologyreview.org', 'www.fao.org', 'www.ijhssi.org', ['journal of ethnic foods'], ['[[gastronomica'], ['gastronomica'], ['poultry science '], ['poultry science'], [' genetics selection evolution '], ['gastronomica'], ['[[journal of heredity'], ['journal of the experimental analysis of behavior']]",15920272,Allow all users (no expiry set),29381,24 February 2008,Steven Walling ,545,1,2008-02-24,2008-02,2008
96,96,Outline of food preparation,https://en.wikipedia.org/wiki/Outline_of_food_preparation,4,0,[],[],1,0,0,2,0,0,1,0.25,0.0,0.5,0.0,0.0,0.25,0,"['www.tescorealfood.com', 'about.com', 'www.fao.org']",3209485,Allow all users (no expiry set),15478,21 November 2005,Go for it! ,455,3,2005-11-21,2005-11,2005
97,97,Provence,https://en.wikipedia.org/wiki/Provence,56,1,"['10.1186/1471-2148-11-69', '21401952', '3068964']",[['bmc evolutionary biology ']],1,0,0,5,0,0,49,0.017857142857142856,0.0,0.08928571428571429,0.017857142857142856,0.0,0.03571428571428571,1,"['kitchen-notebook.blogspot.com', 'nice-cooking.com', 'books.google.com', 'benvengudo.com', 'www.historyofquilts.com', 'www.institut-lumiere.org', ['bmc evolutionary biology ']]",48503,Allow all users (no expiry set),107321,9 April 2002,Pgdudda ,2282,0,2002-04-09,2002-04,2002
98,98,Sauce,https://en.wikipedia.org/wiki/Sauce,16,0,[],[],1,0,0,7,0,0,8,0.0625,0.0,0.4375,0.0,0.0,0.0625,0,"['cooking.nytimes.com', 'uncorneredmarket.com', 'books.google.com', 'books.google.com', 'www.recipetips.com', 'circassianworld.com', 'www.thekitchn.com', 'babel.hathitrust.org']",61937,"Require autoconfirmed or confirmed access (12:50, 11 February 2023)",20404,13 July 2002,Roadrunner ,1920,0,2002-07-13,2002-07,2002
99,99,Delhi,https://en.wikipedia.org/wiki/Delhi,278,4,"['10.1016/j.biocon.2021.109215', None, '10.1093/jue/juab001', '10.2307/604073', None, '25464689', None, None, None, None, None, None]","[['biological conservation'], ['journal of environmental science and engineering '], ['journal of urban ecology'], [' journal of the american oriental society ']]",19,22,0,157,0,2,75,0.0683453237410072,0.07913669064748201,0.564748201438849,0.014388489208633094,0.0,0.1618705035971223,4,"['www.censusindia.gov', 'censusindia.gov', 'censusindia.gov', 'www.archive.india.gov', 'planningcommission.gov', 'www.delhitourism.gov', 'imdpune.gov', 'delhi.gov', 'censusindia.gov', 'city.imd.gov', 'tcpomud.gov', 'mhrd.gov', 'india.gov', 'delhi.gov', 'censusindia.gov', 'censusindia.gov', 'imdpune.gov', 'www.indiapost.gov', 'www.imdpune.gov', 'censusindia.gov', 'pibmumbai.gov', 'unccdcop14india.gov', 'www.indian-handicrafts-suppliers.com', 'www.ndtv.com', 'virsanghvi.com', 'articles.timesofindia.indiatimes.com', 'articles.economictimes.indiatimes.com', 'www.hindustantimes.com', 'cities.expressindia.com', 'indianexpress.com', 'www.hindustantimes.com', 'news.google.com', 'articles.timesofindia.indiatimes.com', 'www.nytimes.com', 'articles.timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'indianexpress.com', 'www.thehindu.com', 'www.cnn.com', 'www.hindustantimes.com', 'timesofindia.indiatimes.com', 'bloomberg.com', 'articles.timesofindia.indiatimes.com', 'www.thehindubusinessline.com', 'www.hindustantimes.com', 'indhistory.com', 'rediff.com', 'delhibarcouncil.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.mapsofindia.com', 'india.blogs.nytimes.com', 'blogs.timesofindia.indiatimes.com', 'indianexpress.com', 'www.ukmediacentre.pwc.com', 'www.indfy.com', 'economictimes.indiatimes.com', 'www.news24.com', 'www.hindustantimes.com', 'mapsofindia.com', 'articles.economictimes.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'economictimes.indiatimes.com', 'www.nytimes.com', 'www.washingtonpost.com', 'www.aboutpalaceonwheels.com', 'in.reuters.com', 'rediff.com', 'www.dailytimes.com', 'delhimetrorail.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.voanews.com', 'books.google.com', 'books.google.com', 'www.indianexpress.com', 'articles.timesofindia.indiatimes.com', 'www.wsj.com', 'timesofindia.indiatimes.com', 'www.reuters.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.news18.com', 'www.apsinghlawyer.com', 'www.nytimes.com', 'kolkatafootballs.com', 'www.hindu.com', 'economictimes.indiatimes.com', 'www.indiatvnews.com', 'outlookindia.com', 'www.mewarindia.com', 'www.economist.com', 'www.espncricinfo.com', 'www.delhimetrorail.com', 'www.terragalleria.com', 'indianexpress.com', 'www.indianexpress.com', 'www.thehindu.com', 'www.hindu.com', 'tribuneindia.com', 'www.nytimes.com', 'www.hindustantimes.com', 'www.washingtonpost.com', 'www.hindu.com', 'www.aipsmedia.com', 'www.economist.com', 'outlookindia.com', 'delhimetrorail.com', 'www.onlineschooladmissions.com', 'www.dailypioneer.com', 'blogs.wsj.com', 'articles.timesofindia.indiatimes.com', 'ndtv.com', 'articles.timesofindia.indiatimes.com', 'www.nytimes.com', 'www.delhimetrorail.com', 'indianexpress.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.niticentral.com', 'economictimes.indiatimes.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.delhimetrorail.com', 'articles.economictimes.indiatimes.com', 'timesofindia.indiatimes.com', 'blogs.wsj.com', 'indlaw.com', 'books.google.com', 'www.hindu.com', 'books.google.com', 'books.google.com', 'www.demographia.com', 'www.india-seminar.com', 'economictimes.indiatimes.com', 'www.indianexpress.com', 'www.dailypioneer.com', 'www.foreignpolicy.com', 'citiesprogramme.com', 'www.hindustantimes.com', 'm.indiatvnews.com', 'www.business-standard.com', 'www.hindu.com', 'books.google.com', 'in.reuters.com', 'books.google.com', 'weatherspark.com', 'timesofindia.indiatimes.com', 'articles.economictimes.indiatimes.com', 'timesofindia.indiatimes.com', 'avalanchepress.com', 'books.google.com', 'airport-delhi.com', 'www.business-standard.com', 'books.google.com', 'economictimes.indiatimes.com', 'books.google.com', 'books.google.com', 'newsfeed.time.com', 'www.hindu.com', 'timesofindia.indiatimes.com', 'www.vidhyasociety.com', 'www.clbuzz.com', 'world.time.com', 'moneycontrol.com', 'ndtv.com', 'www.hindustantimes.com', 'books.google.com', 'books.google.com', 'www.dnaindia.com', 'indianexpress.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'www.weatherbase.com', 'whc.unesco.org', 'www.digital-development-debates.org', 'tourism.org', 'www.afghanistan-analysts.org', 'hdi.globaldatalab.org', 'www.un.org', 'www.worldcat.org', 'www.digital-development-debates.org', 'cseindia.org', 'www.prsindia.org', 'ocasia.org', 'www.cleanairnet.org', 'ocasia.org', 'www.cwgdelhi2010.org', 'whc.unesco.org', 'portal.unesco.org', 'www.undp.org', 'www.downtoearth.org', 'rbidocs.rbi.org', ['biological conservation'], ['journal of environmental science and engineering '], ['journal of urban ecology'], [' journal of the american oriental society ']]",37756,Require autoconfirmed or confirmed access (no expiry set),208265,5 February 2002,Sjc ,12184,16,2002-02-05,2002-02,2002
100,100,Garum,https://en.wikipedia.org/wiki/Garum,39,4,"['10.1093/jhmas/39.4.430', '10.1002/jsfa.1013', '10.1017/s0031182015001651', '6389686', None, '26741568', None, None, None]","[['journal of the history of medicine and allied sciences '], ['journal of the science of food and agriculture'], ['parasitology ']]",4,0,0,12,0,0,19,0.10256410256410256,0.0,0.3076923076923077,0.10256410256410256,0.0,0.20512820512820512,3,"['books.google.com', 'www.timesofisrael.com', 'google.com', 'www.latimes.com', 'books.google.com', 'books.google.com', 'www.salon.com', 'www.haaretz.com', 'books.google.com', 'www.bbc.com', 'books.google.com', 'dsc.discovery.com', 'www.pompeiana.org', 'www.npr.org', 'cooks.aadl.org', 'www.jstor.org', ['journal of the history of medicine and allied sciences '], ['journal of the science of food and agriculture'], ['parasitology ']]",312320,Allow all users (no expiry set),20331,5 September 2003,Ihcoyc ,561,2,2003-09-05,2003-09,2003
101,101,List of English words of Arabic origin,https://en.wikipedia.org/wiki/List_of_English_words_of_Arabic_origin,11,0,[],[],0,0,0,7,0,0,4,0.0,0.0,0.6363636363636364,0.0,0.0,0.0,0,"['baheyeldin.com', 'dict.yulghun.com', 'dict.yulghun.com', '001300-www.al-mostafa.com', 'books.google.com', 'www.m-w.com', 'al-mostafa.com']",574499,Allow all users (no expiry set),31992,3 April 2004,Jengod ,2254,0,2004-04-03,2004-04,2004
102,102,Nice,https://en.wikipedia.org/wiki/Nice,57,3,"['10.1016/0160-7383(79)90095-1', '10.1111/j.1475-4754.1977.tb00189.x', '10.1093/ehr/cxi.433.1018', None, None, None, None, None, None]","[['annals of tourism research '], ['[[archaeometry'], ['the english historical review ']]",2,2,0,15,0,0,35,0.03508771929824561,0.03508771929824561,0.2631578947368421,0.05263157894736842,0.0,0.12280701754385964,3,"['astana.gov', 'www.edinburgh.gov', 'demographia.com', 'www.bestofniceblog.com', 'www.cnn.com', 'www.reuters.com', 'www.startribune.com', 'villeneuveloubethotelreservation.com', 'waybackmachine.com', 'robertwservice.blogspot.com', 'www.france24.com', 'connexionfrance.com', 'www.olympicnice.com', 'www.weather-atlas.com', 'europe-cities.com', 'francemonthly.com', 'www.lejazzophone.com', 'www.musee-terra-amata.org', 'www.nobelprize.org', ['annals of tourism research '], ['[[archaeometry'], ['the english historical review ']]",47088,Allow all users (no expiry set),86947,1 April 2002,WojPob ,4245,8,2002-04-01,2002-04,2002
103,103,Calabria,https://en.wikipedia.org/wiki/Calabria,173,4,"['10.1086/362608', '10.1016/0012-8252(95)00009-7', '10.1021/jf2050075', None, None, '22458691', None, None, None]","[['classical philology'], ['earth-science reviews '], ['j. agric. food chem.']]",6,2,0,64,0,1,96,0.03468208092485549,0.011560693641618497,0.3699421965317919,0.023121387283236993,0.0,0.06936416184971098,3,"['nasa.gov', 'www.burwood.nsw.gov', 'www.intowine.com', 'books.google.com', 'discoveries-in-sicily-and-calabria.blogspot.com', 'www.italyaround.com', 'www.nytimes.com', 'www.madeinsouthitalytoday.com', 'en.italy-holiday.com', 'www.naplesldm.com', 'www.italy24.ilsole24ore.com', 'www.nytimes.com', 'orthochristian.com', 'books.google.com', 'www.timeanddate.com', 'www.panoramitalia.com', 'www.collinsdictionary.com', 'youritaly.com', 'theoi.com', 'www.consorziocipollatropeaigp.com', 'smaf-ltd.com', 'artisanvineyards.com', 'www.italytraveller.com', 'viaggiart.com', 'www.insidersabroad.com', 'bleedingespresso.com', 'www.ethnologue.com', 'www.britannica.com', 'bleedingespresso.com', 'www.youtube.com', 'globalepicurean.com', 'www.deliciousitaly.com', 'vino-con-vista.blogspot.com', 'books.google.com', 'www.freshplaza.com', 'napavalleyregister.com', 'books.google.com', 'www.g-site.com', 'www.amalficoast.com', 'www.greatitalianchefs.com', 'www.italymagazine.com', 'www.dnainfo.com', 'initalytoday.com', 'rabbibarbara.com', 'agronotizie.imagelinenetwork.com', 'www.youtube.com', 'www.youtube.com', 'oliveoilsindia.com', 'www.irishtimes.com', 'www.italy24.ilsole24ore.com', 'www.madeinsouthitalytoday.com', 'www.praiaartresort.com', 'books.google.com', 'www.youtube.com', 'www.givaudan.com', 'eu.greekreporter.com', 'ww1.prweb.com', 'books.google.com', 'www.consorziocipollatropeaigp.com', 'www.britannica.com', 'ourlivesinitaly.com', 'www.youtube.com', 'www.naplesldm.com', 'susanvanallen.wordpress.com', 'highestbridges.com', 'www.railwaypro.com', 'www.olympic.org', 'orthodoxengland.org', 'ftp.fao.org', 'hdi.globaldatalab.org', 'modeoflife.org', 'www.dantemass.org', ['classical philology'], ['earth-science reviews '], ['j. agric. food chem.']]",44772,Allow all users (no expiry set),125691,18 March 2002,62.98.20.244 ,2992,1,2002-03-18,2002-03,2002
104,104,Western India,https://en.wikipedia.org/wiki/Western_India,22,0,[],[],4,3,0,8,0,0,7,0.18181818181818182,0.13636363636363635,0.36363636363636365,0.0,0.0,0.3181818181818182,0,"['www.cia.gov', 'www.gsi.gov', 'www.censusindia.gov', 'books.google.com', 'books.google.com', 'wzccindia.com', 'outlookindia.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.ccsindia.org', 'www.nfhsindia.org', 'www.commonlii.org', 'www.lilaproject.org']",2978812,Allow all users (no expiry set),21496,23 October 2005,2fort5r ,647,5,2005-10-23,2005-10,2005
105,105,Brittany,https://en.wikipedia.org/wiki/Brittany,88,1,"['10.4312/dp.31.8', None, None]",[['documenta praehistorica']],14,0,0,15,0,1,57,0.1590909090909091,0.0,0.17045454545454544,0.011363636363636364,0.0,0.17045454545454544,1,"['books.google.com', 'velo.tourismebretagne.com', 'www.linternaute.com', 'www.megalithes-morbihan.com', 'www.rue89.com', 'www.bretonbikes.com', 'www.agencebretagnepresse.com', 'books.google.com', 'books.google.com', 'www.ifop.com', 'www.festival-interceltique.com', 'emgann.chez.com', 'www.ifop.com', 'www.breizh-amerika.com', 'us.franceguide.com', 'www.ofis-bzh.org', 'www.bretagne-environnement.org', 'www.bretagne-environnement.org', 'www.espace-sciences.org', 'www.espace-sciences.org', 'newgtlds.icann.org', 'www.bretagne-environnement.org', 'bretagne-environnement.org', 'bretagne-environnement.org', 'www.bretagne-environnement.org', 'www.espace-sciences.org', 'www.espace-sciences.org', 'www.prefics.org', 'www.diwanbreizh.org', ['documenta praehistorica']]",38748,Allow all users (no expiry set),127764,11 February 2002,Jeronimo ,3593,5,2002-02-11,2002-02,2002
106,106,Culture of India,https://en.wikipedia.org/wiki/Culture_of_India,204,12,"['10.1111/j.1467-9744.2012.01274.x', '10.1080/15570274.2016.1184437', '10.1038/nature08365', '10.1111/1467-8462.12143', '10.1177/0262728004042760', '10.1093/molbev/msh151', '10.2307/1397540', '10.1080/08949460490274013', '10.1007/s12126-020-09401-x', '10.1093/obo/9780195399318-0071', '10.2307/3250226', '10.2307/2754275', None, None, '19779445', None, None, '15128876', None, None, None, None, None, None, None, None, '2842210', None, None, None, None, None, None, None, None, None]","[['zygon '], ['the review of faith '], ['nature'], ['australian economic review'], ['south asia research'], ['molecular biology and evolution'], ['philosophy east and west '], ['visual anthropology'], ['ageing international '], ['oxford university press '], ['artibus asiae'], ['pacific affairs ']]",19,3,0,75,0,0,95,0.09313725490196079,0.014705882352941176,0.36764705882352944,0.058823529411764705,0.0,0.16666666666666666,12,"['www.fas.usda.gov', 'india.gov', 'www.india.gov', 'www.britannica.com', 'books.google.com', 'www.curiouscook.com', 'www.thehindu.com', 'www.ft.com', 'www.phillipzarrilli.com', 'books.google.com', 'books.google.com', 'books.google.com', 'theflavoursofhistory.com', 'books.google.com', 'www.spectrumcommodities.com', 'books.google.com', 'books.google.com', 'atimes.com', 'www.curiouscook.com', 'www.ibtimes.com', 'www.orissany.com', 'www.hindustantimes.com', 'www.fifa.com', 'bbcvietnamese.com', 'books.google.com', 'books.google.com', 'books.google.com', 'indianpolo.com', 'www.business-standard.com', 'www.meatlessmonday.com', 'books.google.com', 'zawaj.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.ft.com', 'timesofindia.indiatimes.com', 'books.google.com', 'economictimes.indiatimes.com', 'www.indiantelevision.com', 'www.britannica.com', 'books.google.com', 'www.indiapolo.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'www.firstpost.com', 'www.indiantelevision.com', 'ejmas.com', 'www.reuters.com', 'books.google.com', 'indianfoodforever.com', 'www.accessmylibrary.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'www.oup.com', 'books.google.com', 'www.amazon.com', 'spicediary.com', 'www.etymonline.com', 'books.google.com', 'bahai-library.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.iakoweb.com', 'zeenews.india.com', 'books.google.com', 'www.cbsnews.com', 'books.google.com', 'www.icdf.com', 'www.hindu.com', 'www.uniindia.com', 'books.google.com', 'formula1.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.cambridge.org', 'whc.unesco.org', 'whc.unesco.org', 'whc.unesco.org', 'nrn.org', 'whc.unesco.org', 'www.shrm.org', 'whc.unesco.org', 'whc.unesco.org', 'www.cambridge.org', 'www.factsaboutindia.org', 'www.jstor.org', 'www.science.org', 'whc.unesco.org', 'unstats.un.org', 'religioustolerance.org', 'www.cambridge.org', 'sanskritdocuments.org', 'news.bahai.org', ['zygon '], ['the review of faith '], ['nature'], ['australian economic review'], ['south asia research'], ['molecular biology and evolution'], ['philosophy east and west '], ['visual anthropology'], ['ageing international '], ['oxford university press '], ['artibus asiae'], ['pacific affairs ']]",293133,Allow all users (no expiry set),150673,10 August 2003,Mowgli~enwiki ,6371,130,2003-08-10,2003-08,2003
107,107,Paris,https://en.wikipedia.org/wiki/Paris,380,1,"['10.1038/srep02153', '23835429', '3703887']",[['scientific reports']],23,1,0,151,0,5,200,0.060526315789473685,0.002631578947368421,0.3973684210526316,0.002631578947368421,0.0,0.06578947368421052,1,"['travel.state.gov', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'france24.com', 'www.weather-atlas.com', 'parisladefense.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'insidermonkey.com', 'books.google.com', 'books.google.com', 'smithsonian.com', 'books.google.com', 'laposte.com', 'www.forbes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'welections.wordpress.com', 'uk.tourisme93.com', 'books.google.com', 'courrierinternational.com', 'books.google.com', 'www.rolandgarros.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.cnn.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.cnn.com', 'www.forbes.com', 'www.meteofrance.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'olympics.com', 'www.airport-world.com', 'books.google.com', 'books.google.com', 'books.google.com', 'press.parisinfo.com', 'www.usatoday.com', 'www.nytimes.com', 'books.google.com', 'www.afp.com', 'books.google.com', 'french.about.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'www.parisdigest.com', 'books.google.com', 'books.google.com', 'sfcitizen.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.ey.com', 'press.parisinfo.com', 'www.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.com', 'japantoday.com', 'books.google.com', 'books.google.com', 'www.optile.com', 'books.google.com', 'books.google.com', 'courrierinternational.com', 'books.google.com', 'www.tripsavvy.com', 'www.reuters.com', 'www.worldatlas.com', 'www.railwaygazette.com', 'paris.com', 'en.parisinfo.com', 'books.google.com', 'www.britannica.com', 'www.globalwoodmarketsinfo.com', 'www.euronews.com', 'www.britannica.com', 'books.google.com', 'www.cimac.com', 'books.google.com', 'www.tripsavvy.com', 'books.google.com', 'books.google.com', 'www.businessweek.com', 'books.google.com', 'books.google.com', 'books.google.com', 'beatdom.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'articles.timesofindia.indiatimes.com', 'gp-investment-agency.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'about-france.com', 'www.linternaute.com', 'books.google.com', 'www.com', 'books.google.com', 'books.google.com', 'books.google.com', 'french.about.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'iexplore.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.andante.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.google.com', 'www.iied.org', 'wayback.archive-it.org', 'whc.unesco.org', 'franceintheus.org', 'jewishdatabank.org', 'whc.unesco.org', 'whc.unesco.org', 'www.cambridge.org', 'whc.unesco.org', 'www.stif.org', 'www.pewresearch.org', 'wayback.archive-it.org', 'www.oecd-ilibrary.org', 'stats.oecd.org', 'www.metmuseum.org', 'whc.unesco.org', 'www.gutenberg.org', 'www.sciencemuseum.org', 'www.nobelprize.org', 'www.adoremus.org', 'oecd.org', 'www.eib.org', 'wayback.archive-it.org', ['scientific reports']]",22989,Require administrator access (no expiry set),283581,6 November 2001,Zundark ,19327,58,2001-11-06,2001-11,2001
108,108,Malayali,https://en.wikipedia.org/wiki/Malayali,116,1,"['10.33306/mjssh/31', None, None]",[['muallim journal of social sciences and humanities']],3,13,0,49,0,0,51,0.02586206896551724,0.11206896551724138,0.4224137931034483,0.008620689655172414,0.0,0.14655172413793102,1,"['www.pmo.gov', 'www.immi.gov', 'censusindia.gov', 'lsi.gov', 'www.censusindia.gov', 'kerala.gov', 'www.nvtc.gov', 'kerala.gov', 'www.censusindia.gov', 'stats.gov', 'www.cbs.gov', 'abs.gov', 'www.censusindia.gov', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'media.johnwiley.com', 'dances.indobase.com', 'books.google.com', 'www.dnaindia.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', '40days.homestead.com', 'books.google.com', 'keralaliterature.com', 'www.thehindu.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.yourdiscovery.com', 'unreachednewyork.com', 'query.nytimes.com', 'books.google.com', 'timesofindia.indiatimes.com', 'food.ndtv.com', 'books.google.com', 'books.google.com', 'outlookindia.com', 'books.google.com', 'indianexpress.com', 'www.viennamalayaleeassociation.com', 'www.hindu.com', 'www.thehindu.com', 'books.google.com', 'www.business-standard.com', 'nihonkairali.com', 'books.google.com', 'timesofindia.indiatimes.com', 'keral.com', 'www.vegrecipesofindia.com', 'profile.id.com', 'www.britannica.com', 'books.google.com', 'www.dnaindia.com', 'www.malayalamresourcecentre.org', 'www.malayalamresourcecentre.org', 'www.malayalamresourcecentre.org', ['muallim journal of social sciences and humanities']]",1258430,Allow all users (no expiry set),67891,9 December 2004,QuartierLatin1968 ,3554,1,2004-12-09,2004-12,2004
109,109,Mulukhiyah,https://en.wikipedia.org/wiki/Mulukhiyah,20,1,"['10.1080/03670244.1981.9990646', None, None]",[['ecology of food and nutrition ']],0,0,0,15,0,0,4,0.0,0.0,0.75,0.05,0.0,0.05,1,"['books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'baheyeldin.com', 'foodsfromafrica.com', 'www.etymonline.com', 'www.latimes.com', 'taste.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', ['ecology of food and nutrition ']]",4314987,Allow all users (no expiry set),18389,8 March 2006,Mb1000 ,629,2,2006-03-08,2006-03,2006
110,110,Turin,https://en.wikipedia.org/wiki/Turin,89,0,[],[],7,0,0,37,0,0,46,0.07865168539325842,0.0,0.4157303370786517,0.0,0.0,0.07865168539325842,0,"['www.com', 'focus2move.com', 'euromonitor.com', 'www.uefa.com', 'citymayors.com', 'www.com', 'www.ukmediacentre.pwc.com', 'citymayors.com', 'intesasanpaolo.com', 'footballderbies.com', 'edition.cnn.com', 'www.acmilan.com', 'italiantourism.com', 'fifa.com', 'www.nybooks.com', 'www.com', 'www.com', 'moovitapp.com', 'en.archive.uefa.com', 'citymayors.com', 'moovitapp.com', 'www.ukmediacentre.pwc.com', 'www.nittoatpfinals.com', 'www.com', 'www.usatoday.com', 'italianrus.com', 'www.bloomberg.com', 'lumiq.com', 'www.uefa.com', 'www.com', 'www.com', 'www.acmilan.com', 'www.smh.com', 'books.google.com', 'www.smh.com', 'www.com', 'www.archaeolink.com', 'www.centroestero.org', 'www.piemontefeel.org', 'creativecommons.org', 'climaintoscana.altervista.org', 'torinofilmfest.org', 'europe.uli.org', 'en.wikisource.org']",19450529,Allow all users (no expiry set),121921,3 February 2002,Espen ,4021,13,2002-02-03,2002-02,2002
111,111,Florence,https://en.wikipedia.org/wiki/Florence,135,2,"['10.1016/s0304-4181(02)00002-7', '10.2343/geochemj.39.531', None, None, None, None]","[['journal of medieval history '], ['geochemical journal ']]",9,1,0,62,0,2,59,0.06666666666666667,0.007407407407407408,0.45925925925925926,0.014814814814814815,0.0,0.08888888888888889,2,"['trove.nla.gov', 'www.auxologia.com', 'travelandleisure.com', 'travelguide.affordabletours.com', 'www.euromonitor.com', 'lonelyplanet.com', 'www.com', 'www.italyperfect.com', 'moovitapp.com', 'moovitapp.com', 'books.google.com', 'www.florence-on-line.com', 'florenceholidays.com', 'www.com', 'italian.about.com', 'giuniversity.wordpress.com', 'www.com', 'www.ilsole24ore.com', 'britannica.com', 'www.chicagotribune.com', 'books.google.com', 'www.forbes.com', 'www.com', 'hvs.com', 'city-getaway.com', 'studymode.com', 'virtualuffizi.com', 'bachtrack.com', 'edition.cnn.com', 'books.google.com', 'www.travelingintuscany.com', 'www.italy24.ilsole24ore.com', 'europe.travelonline.com', 'www.visitflorence.com', 'www.velonation.com', 'languagemonitor.com', 'euromonitor.com', 'www.smithsonianmag.com', 'www.fosterandpartners.com', 'www.com', 'search.barnesandnoble.com', 'books.google.com', 'www.winepros.com', 'www.auxologia.com', 'florence.world-guides.com', 'tourism-review.com', 'www.pastellists.com', 'tourism-review.com', 'www.time.com', 'search.alexanderstreet.com', 'cntraveller.com', 'ucatholic.com', 'cntraveler.com', 'florenceholidays.com', 'tripleman.com', 'www.economist.com', 'books.google.com', 'www.britannica.com', 'www.weather-atlas.com', 'books.google.com', 'britannica.com', 'dailyhomelist.com', 'brunelleschisdome.com', 'www.tate.org', 'whc.unesco.org', 'gcatholic.org', 'palazzostrozzi.org', 'www.footballhistory.org', 'learner.org', 'library.thinkquest.org', 'catholic-hierarchy.org', 'aacupi.org', ['journal of medieval history '], ['geochemical journal ']]",11525,Allow all users (no expiry set),124941,19 November 2001,Anders Torlind ,5645,9,2001-11-19,2001-11,2001
112,112,Koyilandy,https://en.wikipedia.org/wiki/Koyilandy,38,0,[],[],3,3,0,8,0,0,24,0.07894736842105263,0.07894736842105263,0.21052631578947367,0.0,0.0,0.15789473684210525,0,"['lsgkerala.gov', 'censusindia.gov', 'sec.kerala.gov', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'www.britannica.com', 'www.fallingrain.com', 'www.cartage.org', 'malappuramtourism.org', 'pressacademy.org']",3967460,Allow all users (no expiry set),23655,5 February 2006,Kjrajesh ,612,4,2006-02-05,2006-02,2006
113,113,Japan,https://en.wikipedia.org/wiki/Japan,375,34,"['10.1016/j.imic.2012.04.004', '10.1038/jhg.2012.114', '10.1093/ijl/5.1.1', '10.1017/s0033822200031854', '10.2307/2048846', '10.1080/08865655.2011.686969', '10.1023/a:1008688209052', '10.2307/2539100', '10.1007/978-3-319-02320-5_36-2', '10.1080/08920753.2013.865008', '10.1111/pcn.12428', '10.1016/j.je.2016.12.017', '10.1002/ece3.2070', '10.2307/132115', '10.1007/s12544-017-0255-7', '10.1093/acprof:oso/9780198205890.001.0001', '10.1007/978-3-319-02344-1_36', '10.2753/jes1097-203x270245', '10.2307/987685', '10.1080/1343943x.2018.1459752', '10.3390/rel10060377', '10.1007/978-3-319-20591-5_14', '10.1080/13504630.2018.1499225', '10.1111/j.0022-3840.2005.00123.x', '10.3389/feart.2020.00205', '10.1111/1467-9701.00522', '10.1080/08865655.2011.686972', '10.1177/0920203x16665778', '10.18111/wtobarometereng.2020.18.1.5', '10.1155/2017/4107614', '10.1007/s40844-016-0064-z', None, '23135232', None, None, None, None, None, None, None, None, '27487762', '28716381', '27066244', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, '5623034', '4798153', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None]","[['journal of marine and island cultures'], ['journal of human genetics'], ['international journal of lexicography'], ['[[radiocarbon '], ['the far eastern quarterly'], ['journal of borderlands studies'], ['european journal of law and economics'], ['international security'], ['springer'], ['coastal management'], ['psychiatry and clinical neurosciences'], ['journal of epidemiology'], [' ecology and evolution'], ['journal of japanese studies'], ['european transport research review'], ['oxford university press'], ['springer international publishing '], ['japanese economy'], ['journal of the society of architectural historians'], ['plant production science'], ['religions'], ['proceedings of the international conference on social modeling and simulation'], ['social identities'], ['journal of popular culture'], ['frontiers in earth science'], ['the world economy'], ['journal of borderlands studies'], ['china information'], ['unwto', 'unwto world tourism barometer'], ['journal of energy'], ['evolutionary and institutional economics review']]",60,6,0,89,0,4,182,0.16,0.016,0.23733333333333334,0.09066666666666667,0.0,0.26666666666666666,31,"['www.state.gov', 'www.cia.gov', 'www.state.gov', 'solarsystem.nasa.gov', 'www.sec.gov', 'www.loc.gov', 'www.bloomberg.com', 'books.google.com', 'www.forbes.com', 'www.economist.com', 'www.topuniversities.com', 'www.thejakartapost.com', 'www.bbc.com', 'www.cnn.com', 'www.nytimes.com', 'edition.cnn.com', 'www.usatoday.com', 'gamasutra.com', 'books.google.com', 'apnews.com', 'variety.com', 'www.google.com', 'www.bbc.com', 'japantoday.com', 'japantoday.com', 'money.cnn.com', 'japan-forward.com', 'fortune.com', 'books.google.com', 'www.google.com', 'www.nytimes.com', 'www.wsj.com', 'www.fifa.com', 'www.autosport.com', 'books.google.com', 'www.statsf1.com', 'qz.com', 'www.koreaherald.com', 'www.theatlantic.com', 'www.fiba.com', 'www.space.com', 'www.rethinktokyo.com', 'www.tokyoweekender.com', 'www.smithsonianmag.com', 'www.bbc.com', 'www.aljazeera.com', 'books.google.com', 'fortune.com', 'www.space.com', 'www.cnn.com', 'www.frommers.com', 'www.motogp.com', 'books.google.com', 'www.bbc.com', 'nippon.com', 'www.marketwatch.com', 'books.google.com', 'www.theatlantic.com', 'www.christianitytoday.com', 'www.rugbyworldcup.com', 'www.japanherald.com', 'www.theatlantic.com', 'www.bbc.com', 'japantoday.com', 'www.cnn.com', 'www.timeout.com', 'www.asiarugby.com', 'nippon.com', 'www.economist.com', 'www.neimagazine.com', 'www.bbc.com', 'www.wrc.com', 'thediplomat.com', 'www.google.com', 'www.nytimes.com', 'www.reuters.com', 'www.thrillist.com', 'www.bbc.com', 'www.globalfirepower.com', 'www.livescience.com', 'www.bbc.com', 'www.reuters.com', 'www.theatlantic.com', 'www.vice.com', 'nippon.com', 'www.afcasiancup.com', 'www.statista.com', 'www.ecowatch.com', 'www.fitchratings.com', 'nippon.com', 'fortune.com', 'asia.nikkei.com', 'www.cnn.com', 'statisticstimes.com', 'books.google.com', 'www.mathunion.org', 'www.olympic.org', 'data.worldbank.org', 'whc.unesco.org', 'calisphere.org', 'stats.oecd.org', 'data.uis.unesco.org', 'www.fivb.org', 'data.worldbank.org', 'dataunodc.un.org', 'www.metmuseum.org', 'www.metmuseum.org', 'www3.weforum.org', 'www.oecd.org', 'www.nobelprize.org', 'hdr.undp.org', 'www.fao.org', 'data.imf.org', 'ifr.org', 'www.un.org', 'www.cfr.org', 'www.pbs.org', 'www.oxfordenergy.org', 'reports.weforum.org', 'ncee.org', 'data.worldbank.org', 'uis.unesco.org', 'www.oecd.org', 'www.oecd.org', 'data.worldbank.org', 'www.oecd.org', 'www.un.org', 'www.jstor.org', 'www.imf.org', 'www.oecd-ilibrary.org', 'www.visionofhumanity.org', 'www.oecd.org', 'www.metmuseum.org', 'www.jcie.org', 'www.metmuseum.org', 'www.cfr.org', 'gpseducation.oecd.org', 'dataunodc.un.org', 'databank.worldbank.org', 'gpseducation.oecd.org', 'dataunodc.un.org', 'protocol.un.org', 'reports.weforum.org', 'web-japan.org', 'data.worldbank.org', 'data.worldbank.org', 'data.oecd.org', 'www.japansociety.org', 'collections.dma.org', 'dataunodc.un.org', 'globaldiplomacyindex.lowyinstitute.org', 'www.ramsar.org', 'www.worldshipping.org', 'www.nypl.org', 'data.worldbank.org', ['journal of marine and island cultures'], ['journal of human genetics'], ['international journal of lexicography'], ['[[radiocarbon '], ['the far eastern quarterly'], ['journal of borderlands studies'], ['european journal of law and economics'], ['international security'], ['springer'], ['coastal management'], ['psychiatry and clinical neurosciences'], ['journal of epidemiology'], [' ecology and evolution'], ['journal of japanese studies'], ['european transport research review'], ['oxford university press'], ['springer international publishing '], ['japanese economy'], ['journal of the society of architectural historians'], ['plant production science'], ['religions'], ['proceedings of the international conference on social modeling and simulation'], ['social identities'], ['journal of popular culture'], ['frontiers in earth science'], ['the world economy'], ['journal of borderlands studies'], ['china information'], ['unwto', 'unwto world tourism barometer'], ['journal of energy'], ['evolutionary and institutional economics review']]",15573,Require administrator access (no expiry set),165667,31 October 2001,Alan D ,19010,31,2001-10-31,2001-10,2001
114,114,Manti (food),https://en.wikipedia.org/wiki/Manti_(food),29,1,[],[],1,0,0,18,0,0,9,0.034482758620689655,0.0,0.6206896551724138,0.034482758620689655,0.0,0.06896551724137931,0,"['books.google.com', 'books.google.com', 'www.confucianism.com', 'books.google.com', 'www.confucianism.com', 'vimeo.com', 'books.google.com', 'lulu.com', 'books.google.com', 'www.lezzet.com', 'www.fuchsiadunlop.com', 'www.hurriyetdailynews.com', 'books.google.com', 'books.google.com', 'www.hurriyet.com', '100.naver.com', 'books.google.com', 'vimeo.com', 'www.sras.org']",2827095,Allow all users (no expiry set),21381,3 October 2005,Macrakis ,998,3,2005-10-03,2005-10,2005
115,115,Romania,https://en.wikipedia.org/wiki/Romania,356,5,"['10.1038/news.2011.8', '10.1038/s41467-020-19493-3', '10.1017/s0043887100008091', '10.1093/biosci/bix014', '10.1038/469142a', None, '33293507', None, '28608869', '21228844', None, '7723057', None, '5451287', None]","[['nature '], ['nature communications'], ['transitions world politics '], ['bioscience'], ['nature ']]",42,10,0,87,0,3,210,0.11797752808988764,0.028089887640449437,0.2443820224719101,0.014044943820224719,0.0,0.1601123595505618,5,"['cia.gov', 'www.cia.gov', 'eia.gov', 'www.cia.gov', 'www.msd.gov', 'www.msd.gov', '2009-2017.state.gov', 'permanent.access.gpo.gov', 'www.cia.gov', 'lcweb2.loc.gov', 'www.romania-insider.com', 'uefa.com', 'www.nytimes.com', 'www.economist.com', 'books.google.com', 'romania-insider.com', 'www.romania-insider.com', 'ziare.com', 'www.gourmet-european-recipes.com', 'www.altfg.com', 'www.bbc.com', 'www.newsweek.com', 'www.britishpathe.com', 'uefa.com', 'www.wsj.com', 'romaniatourism.com', 'www.statista.com', 'bloodyelbow.com', 'www.fourfourtwo.com', 'ziare.com', 'www.romania-insider.com', 'fightbreak.com', 'www.festival-cannes.com', 'books.google.com', 'www.spacewar.com', 'www.statista.com', 'www.daviscup.com', 'www.schengenvisainfo.com', 'www.theversed.com', 'romania-insider.com', 'ed-u.com', 'www.rsssf.com', 'atptour.com', 'www.bbc.com', 'www.antiquesandthearts.com', 'ceicdata.com', 'indexmundi.com', 'www.bbc.com', 'fourfourtwo.com', 'topuniversities.com', 'www.romania-central.com', 'uefa.com', 'books.google.com', 'educations.com', 'regard-est.com', 'www.bloomberg.com', 'voanews.com', 'romania-insider.com', 'www.eurosport.com', 'books.google.com', 'romaniaturistica.com', 'tribuna.com', 'www.topendsports.com', 'uefa.com', 'uefa.com', 'www.reuters.com', 'travelmakertours.com', 'www.usatoday.com', 'uefa.com', 'www.gheorghe-zamfir.com', 'unseenromania.com', 'www.romania-insider.com', 'aboutromania.com', 'topuniversities.com', 'www.bbc.com', 'www.ainonline.com', 'onejive.com', 'oxfordscholarship.com', 'www.romania-insider.com', 'flightglobal.com', 'acmilanspot.com', 'www.reuters.com', 'gazette.com', 'www.reuters.com', 'query.nytimes.com', 'romania-insider.com', 'www.olympiandatabase.com', 'fifa.com', 'nytimes.com', 'denisamorariu.wordpress.com', 'english.peopledaily.com', 'www.romania-insider.com', 'www.nytimes.com', 'books.google.com', 'www.usatoday.com', 'www.bucharestherald.com', 'indexmundi.com', 'hdr.undp.org', 'whc.unesco.org', 'www3.weforum.org', 'www.imf.org', 'wayback.archive-it.org', 'earthtrends.wri.org', 'pewforum.org', 'europeanregionofgastronomy.org', 'cnewa.org', 'www.unesco.org', 'www.imf.org', 'inwent.org', 'imf.org', 'www.carnivoreconservation.org', 'nobelprize.org', 'transparency.org', 'www.pewforum.org', 'www.imf.org', 'francophonie.org', 'www1.yadvashem.org', 'www.rferl.org', 'www.wilsoncenter.org', 'datahelpdesk.worldbank.org', 'enescusociety.org', 'data.worldbank.org', 'heritage.org', 'nobelprize.org', 'www.imf.org', 'worldbank.org', 'hdr.undp.org', 'www.carnivoreconservation.org', 'ourworldindata.org', 'hdrstats.undp.org', 'www.pewforum.org', 'web.worldbank.org', 'www.wto.org', 'www.worldheritagesite.org', 'www.mdgmonitor.org', 'fao.org', 'whc.unesco.org', 'www.urbanaudit.org', 'www.doingbusiness.org', ['nature '], ['nature communications'], ['transitions world politics '], ['bioscience'], ['nature ']]",25445,Require administrator access (no expiry set),237975,24 March 2001,Rob Salzman ,16032,20,2001-03-24,2001-03,2001
116,116,Jain vegetarianism,https://en.wikipedia.org/wiki/Jain_vegetarianism,19,1,"['10.15273/jue.v2i2.8146', None, None]",[['journal for undergraduate ethnography']],1,0,0,6,0,0,11,0.05263157894736842,0.0,0.3157894736842105,0.05263157894736842,0.0,0.10526315789473684,1,"['www.hindu.com', 'emirates.com', 'atmadrarma.com', 'hinduonnet.com', 'm.food.ndtv.com', 'food.ndtv.com', 'www.pewresearch.org', ['journal for undergraduate ethnography']]",3587235,Allow all users (no expiry set),20554,1 January 2006,DotShell ,498,4,2006-01-01,2006-01,2006
117,117,Peloponnese,https://en.wikipedia.org/wiki/Peloponnese,60,2,"['10.12681/eadd/8139', '10.11141/ia.34.4', None, None, None, None]","[['didaktorika.gr', 'universite des sciences humaines - strasbourg ii'], ['internet archaeology']]",0,0,0,10,0,0,48,0.0,0.0,0.16666666666666666,0.03333333333333333,0.0,0.03333333333333333,2,"['books.google.com', 'books.google.com', 'books.google.com', 'www.nature.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', ['didaktorika.gr', 'universite des sciences humaines - strasbourg ii'], ['internet archaeology']]",45749,Allow all users (no expiry set),50450,24 March 2002,12.255.158.77 ,1144,3,2002-03-24,2002-03,2002
118,118,Apulia,https://en.wikipedia.org/wiki/Apulia,41,2,[],[],2,0,0,17,0,2,18,0.04878048780487805,0.0,0.4146341463414634,0.04878048780487805,0.0,0.0975609756097561,0,"['www.dopitalianfood.com', 'www.oliveoilsitaly.com', 'books.google.com', 'winetourism.com', 'www.oliveoilemporium.com', 'www.gaypugliapodcast.com', 'books.google.com', 'www.winetourism.com', 'www.lonelyplanet.com', 'www.lonelyplanet.com', 'www.thethinkingtraveller.com', 'books.google.com', 'ethnologue.com', 'www.lucerooliveoil.com', 'ethnologue.com', 'www.artecibo.com', 'www.roughguides.com', 'completamente.org', 'hdi.globaldatalab.org']",44783,Allow all users (no expiry set),36683,18 March 2002,62.98.20.244 ,1564,9,2002-03-18,2002-03,2002
119,119,India,https://en.wikipedia.org/wiki/India,226,11,"['10.1017/s0022050709000400', '10.1016/s2542-5196(18)30261-4', '10.1057/s41271-018-0149-5', '10.2305/iucn.uk.2008.rlts.t9917a13026736.en', '10.2307/2645149', '10.2305/iucn.uk.2004.rlts.t58583a11789937.en', '10.2305/iucn.uk.2004.rlts.t54584a11155448.en', '10.1080/085640032000063977', '10.1017/s0007123409990226', '10.2305/iucn.uk.2008.rlts.t44694a10927987.en', '10.1016/j.jhydrol.2018.10.012', None, '30528905', '30353132', None, None, None, None, None, None, None, None, None, '6358127', None, None, None, None, None, None, None, None, None]","[['journal of economic history'], ['[[the lancet planetary health'], ['[[journal of public health policy'], ['[[the iucn red list of threatened species'], ['[[asian survey'], [' [[the iucn red list of threatened species', ' [[iucn'], ['[[the iucn red list of threatened species', '[[iucn'], ['south asia'], ['[[british journal of political science'], ['[[the iucn red list of threatened species'], ['[[journal of hydrology']]",27,20,0,134,0,3,31,0.11946902654867257,0.08849557522123894,0.5929203539823009,0.048672566371681415,0.0,0.25663716814159293,11,"['www.uscirf.gov', 'www.legislative.gov', 'censusindia.gov', 'www.itis.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'dashboard.udiseplus.gov', 'zsi.gov', 'www.censusindia.gov', 'lsi.gov', 'utki.gov', 'rajbhasha.gov', 'www.investindia.gov', 'www.studyinindia.gov', 'www.censusindia.gov', 'www.cia.gov', 'india.gov', 'www.ers.usda.gov', 'india.gov', 'www.indiabudget.gov', 'books.google.com', 'wap.business-standard.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.financialexpress.com', 'books.google.com', 'festivals.indobase.com', 'www.thehindu.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'books.google.com', 'dawn.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'www.wtatennis.com', 'books.google.com', 'www.tribuneindia.com', 'www.thehindu.com', 'hindustantimes.com', 'www.ndtv.com', 'www.news18.com', 'books.google.com', 'www.thehindubusinessline.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.ethnologue.com', 'economictimes.indiatimes.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.britannica.com', 'books.google.com', 'foreignpolicy.com', 'books.google.com', 'www.oed.com', 'books.google.com', 'books.google.com', 'foreignpolicy.com', 'books.google.com', 'www.bbc.com', 'books.google.com', 'www.bbc.com', 'www.financialexpress.com', 'www.thehindubusinessline.com', 'timesofindia.indiatimes.com', 'www.tribuneindia.com', 'www.chessvibes.com', 'indianexpress.com', 'sify.com', 'books.google.com', 'books.google.com', 'books.google.com', 'm.timesofindia.com', 'books.google.com', 'books.google.com', 'articles.economictimes.indiatimes.com', 'books.google.com', 'books.google.com', 'm.timesofindia.com', 'books.google.com', 'books.google.com', 'books.google.com', 'economictimes.indiatimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.deccanherald.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'www.nationalheraldindia.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.thehindu.com', 'www.vox.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'differding.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'timesnownews.com', 'books.google.com', 'books.google.com', 'books.google.com', 'm.timesofindia.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'indianexpress.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'deccanherald.com', 'www.skysports.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www2.deloitte.com', 'www.thehindu.com', 'books.google.com', 'www.sportskeeda.com', 'www.hindu.com', 'books.google.com', 'www.hindu.com', 'www.nation.com', 'books.google.com', 'archive.ethnologue.com', 'books.google.com', 'www.dnaindia.com', 'hdr.undp.org', 'whc.unesco.org', 'www.worldbank.org', 'research.amnh.org', 'research.amnh.org', 'www.americasquarterly.org', 'data.worldbank.org', 'www.imf.org', 'www.ibef.org', 'data.worldbank.org', 'siteresources.worldbank.org', 'www.iucn.org', 'data.worldbank.org', 'www.clgf.org', 'www.iea.org', 'www.climatelinks.org', 'www.bangladeshsociology.org', 'www.unenvironment.org', 'www.globalslaveryindex.org', 'www.ilo.org', 'samaj.revues.org', 'www.biodiversitya-z.org', 'data.worldbank.org', 'imf.org', 'data.worldbank.org', 'transparency.org', 'www.worldbank.org', ['journal of economic history'], ['[[the lancet planetary health'], ['[[journal of public health policy'], ['[[the iucn red list of threatened species'], ['[[asian survey'], [' [[the iucn red list of threatened species', ' [[iucn'], ['[[the iucn red list of threatened species', '[[iucn'], ['south asia'], ['[[british journal of political science'], ['[[the iucn red list of threatened species'], ['[[journal of hydrology']]",14533,Require administrator access (no expiry set),303043,26 October 2001,Corvus13 ,26714,54,2001-10-26,2001-10,2001
120,120,Druze,https://en.wikipedia.org/wiki/Druze,305,14,"['10.1038/nature09103', '10.1525/jps.2000.29.4.02p00787', '10.1111/j.1478-1913.1977.tb03313.x', '10.1179/peq.1988.120.1.26', '10.1016/j.cell.2020.04.024', '10.1126/science.1116815', '10.1002/humu.20077', '10.1371/journal.pone.0002105', '10.1080/0142569900110406', '10.1038/srep35837', '10.2307/605981', '10.1038/srep14484', '10.1080/1369183032000170222', '10.2307/595974', '20531471', None, None, None, '32470400', '16151010', '15300852', '18461126', None, '27848937', None, '26434580', None, None, None, None, None, None, None, None, None, '2324201', None, '5111078', None, '4593049', None, None]","[['nature '], [' journal of palestine studies '], ['muslim world '], ['palestine exploration quarterly'], [' cell '], ['[[science '], ['human mutation '], ['plos one'], [' british journal of sociology of education '], ['scientific reports '], ['journal of the american oriental society'], ['scientific reports'], ['journal of ethnic and migration studies '], ['[[journal of the american oriental society']]",24,7,0,73,0,0,187,0.07868852459016394,0.022950819672131147,0.23934426229508196,0.04590163934426229,0.0,0.14754098360655737,14,"['www1.cbs.gov', '2001-2009.state.gov', 'www.cbs.gov', 'www.abs.gov', 'www1.cbs.gov', 'www.cbs.gov', '2001-2009.state.gov', 'books.google.com', 'books.google.com', 'www.druze.com', 'www.arabamerica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.al-monitor.com', 'www.arabamerica.com', 'books.google.com', 'www.druzesect.com', 'books.google.com', 'www.al-amama.com', 'books.google.com', 'www.economist.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'www.infoplease.com', 'www.syrianhistory.com', 'books.google.com', 'www.sciencedaily.com', 'api.nationalgeographic.com', 'books.google.com', 'books.google.com', 'www.israelnationalnews.com', 'www.britannica.com', 'lexicorient.com', 'tjgorton.wordpress.com', 'books.google.com', 'dictionary.reference.com', 'books.google.com', 'books.google.com', 'english.al-akhbar.com', 'books.google.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'www.cbsnews.com', 'books.google.com', 'www.al-amama.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.middle-east-online.com', 'books.google.com', 'books.google.com', 'www.tabletmag.com', 'books.google.com', 'www.haaretz.com', 'books.google.com', 'thearabweekly.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.latimes.com', 'books.google.com', 'books.google.com', 'www.dailystar.com', 'thestar.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'books.google.com', 'www.al-amama.com', 'books.google.com', 'www.reuters.com', 'www.juf.org', 'books.openedition.org', 'www.eial.org', 'www.idi.org', 'www.druzestudies.org', 'www.iranicaonline.org', 'www.jewishvirtuallibrary.org', 'www.theisraelproject.org', 'weekly.ahram.org', 'www.druzeheritage.org', 'www.refworld.org', 'druzestudies.org', 'www.commentary.org', 'www.internal-displacement.org', 'www.juf.org', 'www.pewforum.org', 'www.druze.org', 'www.sacredtribesjournal.org', 'www.unaids.org', 'www.sacredtribesjournal.org', 'meib.org', 'www.washingtoninstitute.org', 'www.jewishvirtuallibrary.org', 'druze.org', ['nature '], [' journal of palestine studies '], ['muslim world '], ['palestine exploration quarterly'], [' cell '], ['[[science '], ['human mutation '], ['plos one'], [' british journal of sociology of education '], ['scientific reports '], ['journal of the american oriental society'], ['scientific reports'], ['journal of ethnic and migration studies '], ['[[journal of the american oriental society']]",8632,Allow all users (no expiry set),190103,10 October 2001,RK ,4790,19,2001-10-10,2001-10,2001
121,121,Hispanic America,https://en.wikipedia.org/wiki/Hispanic_America,34,4,"['10.1353/hub.2004.0058', None, '10.1093/socrel/srx030', '10.1086/303004', '15754971', '17573655', None, '10873790', None, None, None, '1287189']","[['human biology'], ['genetics and molecular research'], ['sociology of religion'], [' [[the american journal of human genetics']]",9,3,0,6,0,0,12,0.2647058823529412,0.08823529411764706,0.17647058823529413,0.11764705882352941,0.0,0.47058823529411764,4,"['www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'glaniad.com', 'www.crwflags.com', '1stclassargentina.com', 'andesceltig.com', 'patagonline.com', 'www.thefreedictionary.com', 'www.pewforum.org', 'data.worldbank.org', 'www.kacike.org', 'www.pewforum.org', 'data.worldbank.org', 'www.imf.org', 'www.kacike.org', 'argbrit.org', 'www.pewforum.org', ['human biology'], ['genetics and molecular research'], ['sociology of religion'], [' [[the american journal of human genetics']]",452104,Allow all users (no expiry set),47108,2 February 2004,JeLuF ,776,1,2004-02-02,2004-02,2004
122,122,Lesbos,https://en.wikipedia.org/wiki/Lesbos,32,0,[],[],4,1,0,12,0,1,14,0.125,0.03125,0.375,0.0,0.0,0.15625,0,"['dossier.ogp.noaa.gov', 'www.nbcnews.com', 'www.itsaboutgreece.com', 'www.dictionary.com', 'www.nytimes.com', 'greekcitytimes.com', 'www.gamesradar.com', 'www.nationalgeographic.com', 'drive.google.com', 'www.demetrimusic.com', 'www.nationalgeographic.com', 'www.washingtonpost.com', 'greekreporter.com', 'www.wmf.org', 'art.thewalters.org', 'www.globalgeopark.org', 'www.unesco.org']",2633994,Allow all users (no expiry set),40274,7 September 2005,Darwinek ,1936,3,2005-09-07,2005-09,2005
123,123,Frog legs,https://en.wikipedia.org/wiki/Frog_legs,41,0,[],[],4,0,0,30,0,1,6,0.0975609756097561,0.0,0.7317073170731707,0.0,0.0,0.0975609756097561,0,"['www.goodindonesianfood.com', 'books.google.com', 'www.jpnn.com', 'www.villagevoice.com', 'www.exoticmeatsandmore.com', 'www.allmychefs.com', 'nutritiondata.self.com', 'www.lifeinitaly.com', 'www.listsofnote.com', 'konsultasisyariah-akhowatkpii.blogspot.com', 'books.google.com', 'majalah.tempointeraktif.com', 'books.google.com', 'books.google.com', 'books.google.com', 'abcnews.go.com', 'unvegan.com', 'books.google.com', 'books.google.com', 'www.vecer.com', 'books.google.com', 'books.google.com', 'books.google.com', 'issuu.com', 'www.savethefrogs.com', 'books.google.com', 'www.chow.com', 'flavorwire.com', 'www.foodbeast.com', 'issuu.com', 'defenders.org', 'npr.org', 'www.danwei.org', 'eattheinvaders.org']",543812,Allow all users (no expiry set),26807,22 March 2004,203.101.38.241 ,892,2,2004-03-22,2004-03,2004
124,124,Rhodes,https://en.wikipedia.org/wiki/Rhodes,84,2,"['10.1007/s11598-006-9014-9', '10.1023/a:1009706415417', None, None, None, None]","[[' human evolution '], ['[[journal of seismology']]",4,2,0,11,0,0,65,0.047619047619047616,0.023809523809523808,0.13095238095238096,0.023809523809523808,0.0,0.09523809523809523,2,"['www.mfa.gov', 'ftp.atdd.noaa.gov', 'catholicchurchrhodes.com', 'www.milliyet.com', 'www.batitrakya.4mg.com', 'www.britannica.com', 'www.greeka.com', 'books.google.com', 'www.discover-rhodes.com', 'books.google.com', 'www.weather-atlas.com', 'dadfetured.blogspot.com', 'boat-cruises-trips.com', 'jewishvirtuallibrary.org', 'jewishvirtuallibrary.org', 'www.duhaime.org', 'constitution.org', [' human evolution '], ['[[journal of seismology']]",26773183,Allow all users (no expiry set),88178,9 March 2002,Pgdudda ,1835,4,2002-03-09,2002-03,2002
125,125,Nepal,https://en.wikipedia.org/wiki/Nepal,366,23,"['10.2307/2760015', '10.1111/j.1365-2117.2006.00305.x', '10.1038/s41467-020-19493-3', '10.1111/j.1365-246x.2004.02038.x', None, '10.3126/on.v6i1.1657', '10.1016/j.jseaes.2005.10.016', '10.3126/dsaj.v12i0.22176', '10.3126/dsaj.v1i0.284', '10.1016/s1367-9120(99)00034-6', '10.1016/j.jenvman.2014.07.047', '10.1029/94jb00714', '10.1186/s13002-017-0148-9', '10.3126/rnjds.v1i2.22425', '10.3126/nccj.v4i1.24741', '10.2307/2645740', '10.1111/j.1365-246x.2004.02180.x', '10.1016/j.earscirev.2005.07.005', '10.1017/s0041977x00002007', '10.1017/cbo9780511807251.008', '10.1038/jhg.2012.8', '10.3126/jps.v18i0.20439', None, None, '33293507', None, None, None, None, None, None, None, '25181944', None, '28356115', None, None, None, None, None, None, None, '22437208', None, None, None, '7723057', None, 'org/abstract/cba/371633', None, None, None, None, None, None, None, '5372287', None, None, None, None, None, None, None, None, None]","[['pacific affairs '], ['basin research '], ['nature communications '], ['geophys. j. int. '], ['acta botanica yunnanica '], ['our nature '], ['journal of asian earth sciences '], ['dhaulagiri journal of sociology and anthropology'], ['[[dhaulagiri journal of sociology and anthropology'], ['journal of asian earth sciences '], ['journal of environmental management '], ['[[journal of geophysical research'], ['journal of ethnobiology and ethnomedicine '], ['research nepal journal of development studies'], ['ncc journal'], ['[[asian survey'], ['geophys. j. int. '], ['earth-science reviews'], ['bulletin of the school of oriental and african studies'], ['games of no chance ', '[[msri publications'], ['journal of human genetics'], ['[[journal of political science']]",71,23,0,181,0,1,67,0.19398907103825136,0.06284153005464481,0.49453551912568305,0.06284153005464481,0.0,0.319672131147541,22,"['nkp.gov', 'mofa.gov', 'mofa.gov', 'nhrc.gov', 'nta.gov', 'www.cia.gov', 'www.lawcommission.gov', 'www.cia.gov', 'pubs.usgs.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'mohp.gov', 'www.cia.gov', 'np.usembassy.gov', 'cbs.gov', 'mea.gov', 'mofa.gov', 'mofa.gov', 'www.loc.gov', 'tourism.gov', 'moe.gov', 'cbs.gov', 'nepalitimes.com', 'books.google.com', 'english.onlinekhabar.com', 'kathmandupost.com', 'encarta.msn.com', 'nepalnature.com', 'thehimalayantimes.com', 'en.setopati.com', 'admin.myrepublica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'thehimalayantimes.com', 'www.britannica.com', 'kathmandupost.com', 'kathmandupost.com', 'books.google.com', 'narimag.com', 'www.beliefnet.com', 'www.fifa.com', 'kathmandupost.com', 'www.xinhuanet.com', 'archive.nepalitimes.com', 'kathmandupost.ekantipur.com', 'thehimalayantimes.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.espncricinfo.com', 'kathmandupost.com', 'thehimalayantimes.com', 'nepalitimes.com', 'books.google.com', 'thehimalayantimes.com', 'timesofindia.indiatimes.com', 'books.google.com', 'in.reuters.com', 'www.nytimes.com', 'thehimalayantimes.com', 'thehimalayantimes.com', 'www.latimes.com', 'kathmandupost.com', 'www.icc-cricket.com', 'myrepublica.nagariknetwork.com', 'books.google.com', 'kathmandupost.com', 'www.britannica.com', 'www.nepalitimes.com', 'thehimalayantimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'thehimalayantimes.com', 'books.google.com', 'www.kpmalla.com', 'books.google.com', 'thehimalayantimes.com', 'myrepublica.nagariknetwork.com', 'www.aljazeera.com', 'myrepublica.nagariknetwork.com', 'books.google.com', 'myrepublica.nagariknetwork.com', 'kathmandupost.com', 'thehimalayantimes.com', 'books.google.com', 'myrepublica.nagariknetwork.com', 'kathmandupost.com', 'www.latimes.com', 'www.espncricinfo.com', 'kathmandupost.com', 'books.google.com', 'thehimalayantimes.com', 'www.hindu.com', 'kathmandupost.com', 'kathmandupost.com', 'kathmandupost.com', 'thehimalayantimes.com', 'thehimalayantimes.com', 'thehimalayantimes.com', 'books.google.com', 'myrepublica.nagariknetwork.com', 'thediplomat.com', 'kathmandupost.com', 'books.google.com', 'www.nepalitimes.com', 'www.britannica.com', 'english.onlinekhabar.com', 'www.icc-cricket.com', 'kathmandupost.com', 'thediplomat.com', 'books.google.com', 'books.google.com', 'thehimalayantimes.com', 'thehimalayantimes.com', 'kathmandupost.com', 'thehimalayantimes.com', 'myrepublica.nagariknetwork.com', 'thehimalayantimes.com', 'myrepublica.nagariknetwork.com', 'www.espncricinfo.com', 'thehimalayantimes.com', 'books.google.com', 'royalnepal.synthasite.com', 'books.google.com', 'kathmandupost.com', 'books.google.com', 'www.aljazeera.com', 'books.google.com', 'thehimalayantimes.com', 'edusanjal.com', 'books.google.com', 'books.google.com', 'www.bbc.com', 'www.ktm2day.com', 'books.google.com', 'www.aljazeera.com', 'myrepublica.nagariknetwork.com', 'www.reuters.com', 'www.onlinekhabar.com', 'kathmandupost.ekantipur.com', 'kathmandupost.ekantipur.com', 'books.google.com', 'books.google.com', 'www.economist.com', 'books.google.com', 'kathmandupost.com', 'www.nytimes.com', 'www.statista.com', 'www.nepalitimes.com', 'thehimalayantimes.com', 'www.espncricinfo.com', 'books.google.com', 'www.cnn.com', 'www.nepalitimes.com', 'myrepublica.nagariknetwork.com', 'thehimalayantimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.washingtonpost.com', 'www.nepalitimes.com', 'thehimalayantimes.com', 'www.aljazeera.com', 'thehimalayantimes.com', 'kathmandupost.com', 'kathmandupost.com', 'thehimalayantimes.com', 'thehimalayantimes.com', 'kathmandupost.com', 'www.hindustantimes.com', 'myrepublica.nagariknetwork.com', 'www.aljazeera.com', 'www.lexico.com', 'archive.nepalitimes.com', 'cricketarchive.com', 'thehimalayantimes.com', 'books.google.com', 'kathmandupost.com', 'edition.cnn.com', 'books.google.com', 'thehimalayantimes.com', 'thehimalayantimes.com', 'myrepublica.nagariknetwork.com', 'thediplomat.com', 'thehimalayantimes.com', 'myrepublica.nagariknetwork.com', 'www.nepalitimes.com', 'www.fifa.com', 'www.bbc.com', 'www.infoplease.com', 'kathmandupost.com', 'books.google.com', 'www.sportskeeda.com', 'kathmandupost.com', 'kathmandupost.com', 'books.google.com', 'myrepublica.nagariknetwork.com', 'books.google.com', 'books.google.com', 'thehimalayantimes.com', 'books.google.com', 'thehimalayantimes.com', 'ourworldindata.org', 'www.mhtf.org', 'therisingnepal.org', 'ihl-databases.icrc.org', 'birdlifenepal.org', 'nepal.unfpa.org', 'therisingnepal.org', 'www.globalslaveryindex.org', 'www.adb.org', 'www.wto.org', 'data.worldbank.org', 'www.greenleft.org', 'nc.iucnredlist.org', 'projects.worldbank.org', 'www.unhcr.org', 'www.iucn.org', 'data.worldbank.org', 'therisingnepal.org', 'www.worldbank.org', 'unesdoc.unesco.org', 'hdr.undp.org', 'data.worldbank.org', 'nc.iucnredlist.org', 'reporting.unhcr.org', 'nepal.unfpa.org', 'therisingnepal.org', 'hdrstats.undp.org', 'www.therisingnepal.org', 'www.saferworld.org', 'niss.org', 'peacekeeping.un.org', 'data.worldbank.org', 'data.worldbank.org', 'www.unicef.org', 'therisingnepal.org', 'data.worldbank.org', 'therisingnepal.org', 'www.pewforum.org', 'data.worldbank.org', 'data.worldbank.org', 'www.worldbank.org', 'www.ramsar.org', 'data.worldbank.org', 'www.imf.org', 'www.wwfnepal.org', 'www.imf.org', 'therisingnepal.org', 'www.thenewhumanitarian.org', 'www.unhcr.org', 'whc.unesco.org', 'www.unicef.org', 'www.ilo.org', 'www.imf.org', 'www.wwfnepal.org', 'data.worldbank.org', 'asiafoundation.org', 'www.unhcr.org', 'sari-energy.org', 'www.iucn.org', 'www.worldbank.org', 'data.worldbank.org', 'reporting.unhcr.org', 'csw.org', 'cdm15738.contentdm.oclc.org', 'data.worldbank.org', 'www.internal-displacement.org', 'uis.unesco.org', 'therisingnepal.org', 'visionofhumanity.org', 'asiafoundation.org', 'www.deathpenalty.org', ['pacific affairs '], ['basin research '], ['nature communications '], ['geophys. j. int. '], ['acta botanica yunnanica '], ['our nature '], ['journal of asian earth sciences '], ['dhaulagiri journal of sociology and anthropology'], ['[[dhaulagiri journal of sociology and anthropology'], ['journal of asian earth sciences '], ['journal of environmental management '], ['[[journal of geophysical research'], ['journal of ethnobiology and ethnomedicine '], ['research nepal journal of development studies'], ['ncc journal'], ['[[asian survey'], ['geophys. j. int. '], ['earth-science reviews'], ['bulletin of the school of oriental and african studies'], ['games of no chance ', '[[msri publications'], ['journal of human genetics'], ['[[journal of political science']]",171166,Require administrator access (no expiry set),233655,25 May 2001,KoyaanisQatsi ,8638,8,2001-05-25,2001-05,2001
126,126,Italy,https://en.wikipedia.org/wiki/Italy,631,12,"['10.2307/367499', '10.7551/mitpress/9780262019613.001.0001', '10.1057/9781137008695_19', '10.1038/ejcn.2017.58', '10.1051/ocl.2000.0077', '10.1038/sdata.2018.214', '10.1016/j.jhevol.2011.11.009', '10.1002/wow3.54', '10.2307/1170959', '10.1038/s41467-020-19493-3', '10.5195/jwsr.2006.369', '10.1017/s0033822200040534', None, None, None, '28488692', None, '30375988', '22189428', None, None, '33293507', None, None, None, None, None, None, None, '6207062', None, None, None, '7723057', None, None]","[['history of education quarterly '], ['mit press '], ['palgrave macmillan '], ['european journal of clinical nutrition '], ['oléagineux'], ['scientific data '], [' journal of human evolution '], ['world of work report'], ['social science history '], ['nature communications'], ['journal of world-systems research '], ['radiocarbon ']]",60,13,0,167,0,7,377,0.09508716323296355,0.020602218700475437,0.26465927099841524,0.01901743264659271,0.0,0.1347068145800317,12,"['www.mit.gov', 'factfinder.census.gov', 'www.fco.gov', 'www.sicurezzanazionale.gov', 'www.export.gov', 'www.mite.gov', 'www.salute.gov', 'www.censusdata.abs.gov', 'unmig.sviluppoeconomico.gov', 'www.fco.gov', 'www.cia.gov', 'www.cia.gov', 'www.loc.gov', 'birn.eu.com', 'www.france24.com', 'books.google.com', 'it.yourtripagent.com', 'books.google.com', 'stanzedicinema.com', 'archive.nytimes.com', 'www.sorrisi.com', 'www.economist.com', 'www.britannica.com', 'nriinternet.com', 'articles.sun-sentinel.com', 'books.google.com', 'www.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'languagemonitor.com', 'www.esctoday.com', 'www.boston.com', 'www.history.com', 'dot.com', 'www.bbc.com', 'www.britannica.com', 'ilsole24ore.com', 'nytimes.com', 'www.hotelsclick.com', 'nytimes.com', 'airwaysmag.com', 'books.google.com', 'books.google.com', 'www.shanghairanking.com', 'bestofsicily.com', 'worldpopulationreview.com', 'inmamaskitchen.com', 'books.google.com', 'www.economist.com', 'britannica.com', 'books.google.com', 'books.google.com', 'www.faretennis.com', 'www.ft.com', 'www.oldcalculatormuseum.com', 'www.com', 'www.britannica.com', 'books.google.com', 'www.eni.com', 'books.google.com', 'nationmaster.com', 'italytravel.com', 'adnkronos.com', 'books.google.com', 'adnkronos.com', 'encyclopedia.com', 'www.huffingtonpost.com', 'books.google.com', 'www.britannica.com', 'giornalevinocibo.com', 'www.vogue.com', 'fifa.com', 'www.nytimes.com', 'www.viaggiarenews.com', 'acea.thisconnect.com', 'books.google.com', 'www.economist.com', 'www.nytimes.com', 'www.britannica.com', 'www.wiley.com', 'books.google.com', 'italoamericano.com', 'www.oldcalculatormuseum.com', 'www.com', 'www.timescolonist.com', 'www.antimafiaduemila.com', 'britannica.com', 'adnkronos.com', 'books.google.com', 'www.enel.com', 'www.oldcalculatormuseum.com', 'www.moviemaker.com', 'finance.yahoo.com', 'www.economist.com', 'books.google.com', 'www.bbc.com', 'f1ingenerale.com', 'www.cnbc.com', 'books.google.com', 'epicurean.com', 'www.dw.com', 'www.britannica.com', 'www.hellenicshippingnews.com', 'www.hollywoodreporter.com', 'books.google.com', 'www.dw.com', 'dev.prenhall.com', 'brandfinance.com', 'www.statista.com', 'britannica.com', 'indigoguide.com', 'www.travelpulse.com', 'photius.com', 'www.nytimes.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'art-and-archaeology.com', 'books.google.com', 'www.britannica.com', 'italytravel.com', 'www.bbc.com', 'books.google.com', 'www.nytimes.com', 'www.frieze.com', 'www.uciprotour.com', 'www.italy24.ilsole24ore.com', 'books.google.com', 'www.reuters.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.leithart.com', 'books.google.com', 'www.google.com', 'criterion.com', 'www.britannica.com', 'time.com', 'jakubmarian.com', 'rusticocooking.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.museoauto.com', 'www.harrisinteractive.com', 'www.history.com', 'www.homolaicus.com', 'uk.reuters.com', 'www.britannica.com', 'filmreference.com', 'sallybernstein.com', 'www.solarserver.com', 'www.worldatlas.com', 'catalogue-lumiere.com', 'www.cnbc.com', 'wardsauto.com', 'www.ingentaconnect.com', 'www.turismo-oggi.com', 'www.photius.com', 'www.powerhousemuseum.com', 'www.nationsencyclopedia.com', 'dev.prenhall.com', '(8.com', 'www.ilsole24ore.com', 'www.britannica.com', 'ngm.nationalgeographic.com', 'www.adnkronos.com', 'books.google.com', 'edition.cnn.com', 'economicreconstruction.com', 'ethnologue.com', 'italytravel.com', 'www.reuters.com', 'travel.cnn.com', 'rogerebert.suntimes.com', 'www.allempires.com', 'www.amusingplanet.com', 'italytravel.com', 'www.britannica.com', 'library.thinkquest.org', 'whc.unesco.org', 'www.imf.org', 'www.oecd.org', 'www.crvp.org', 'mdgs.un.org', 'databank.worldbank.org', 'amshq.org', 'www.wttc.org', 'www.un.org', 'data.worldbank.org', 'web.worldbank.org', 'stats.oecd.org', 'www.unesco.org', 'nobelprize.org', 'unterm.un.org', 'www.operaamerica.org', 'www.justitaly.org', 'www.pewforum.org', 'history-world.org', 'data.worldbank.org', 'martinprosperity.org', 'www.fastionline.org', 'www.newadvent.org', 'whc.unesco.org', 'beyondforeignness.org', 'www.nrdc.org', 'www.imf.org', 'www.wwindea.org', 'new.sis-statistica.org', 'www.unesco.org', 'unstats.un.org', 'library.thinkquest.org', 'hdr.undp.org', 'www.world-nuclear.org', 'ourworldindata.org', 'hdr.undp.org', 'www.eurojewcong.org', 'biotaxa.org', 'flpdifesa.org', 'www.dartmouthapologia.org', 'www.chiesavaldese.org', 'www.iotf.org', 'whc.unesco.org', 'www.eoearth.org', 'www.globalwitness.org', 'www.justitaly.org', 'www.oikoumene.org', 'unesco.org', 'metmuseum.org', 'www.oecd.org', 'www.imf.org', 'openknowledge.worldbank.org', 'www.unesco.org', 'www.eurobserv-er.org', 'www.oecd.org', 'databank.worldbank.org', 'www.justitaly.org', 'whc.unesco.org', 'www.justitaly.org', ['history of education quarterly '], ['mit press '], ['palgrave macmillan '], ['european journal of clinical nutrition '], ['oléagineux'], ['scientific data '], [' journal of human evolution '], ['world of work report'], ['social science history '], ['nature communications'], ['journal of world-systems research '], ['radiocarbon ']]",14532,Require administrator access (no expiry set),394172,12 November 2001,Zundark ,18140,109,2001-11-12,2001-11,2001
127,127,Kashk,https://en.wikipedia.org/wiki/Kashk,26,3,"['10.1080/10942912.2018.1466323', '10.1525/gfc.2016.16.4.97', '10.1017/s0022029911000872', None, None, '23171586', None, None, None]","[['international journal of food properties '], ['gastronomica'], ['journal of dairy research ']]",5,0,0,7,0,2,9,0.19230769230769232,0.0,0.2692307692307692,0.11538461538461539,0.0,0.3076923076923077,3,"['jewishstandard.timesofisrael.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'maxima-library.org', 'www.fao.org', 'www.cshd.org', 'www.cshd.org', 'maxima-library.org', ['international journal of food properties '], ['gastronomica'], ['journal of dairy research ']]",3024049,Allow all users (no expiry set),21823,29 October 2005,203.7.227.41 ,397,0,2005-10-29,2005-10,2005
128,128,Indian people,https://en.wikipedia.org/wiki/Indian_people,155,9,"['10.1016/j.ajhg.2013.07.006', '10.1111/j.1475-4754.2008.00454.x', '10.2307/1397540', '10.1016/j.ajhg.2011.11.010', '10.1038/457945a', '10.2307/2053980', '10.2307/2754275', '23932107', None, None, '22152676', '19238684', None, None, '3769933', None, None, '3234374', None, None, None]","[['the american journal of human genetics '], ['archaeometry '], ['philosophy east and west '], ['the american journal of human genetics '], ['nature ', 'nature.com '], [' the journal of asian studies'], ['pacific affairs ']]",14,23,0,37,0,0,72,0.09032258064516129,0.14838709677419354,0.23870967741935484,0.05806451612903226,0.0,0.2967741935483871,7,"['stats.gov', 'pmr.penerangan.gov', 'www.statistics.gov', 'www.statistics.gov', 'www.indembkathmandu.gov', 'www.nationalarchives.gov', 'www.dhs.gov', 'www.uscirf.gov', 'www.dhs.gov', 'moia.gov', 'www.censusindia.gov', 'factfinder.census.gov', 'indembassyisrael.gov', 'www.dhs.gov', 'www.uscirf.gov', 'censusindia.gov', 'mea.gov', 'www.ons.gov', 'www.censusindia.gov', 'www.nationalarchives.gov', 'www.nptd.gov', 'www.dhs.gov', 'www.statssa.gov', 'books.google.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.jerseycityindependent.com', 'bbcvietnamese.com', 'a.harappa.com', 'books.google.com', 'repeatingislands.com', 'books.google.com', 'www.parisschoolofeconomics.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.oup.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'yourarticlelibrary.com', 'gulfnews.com', 'www.sportspundit.com', 'www.milligazette.com', 'tribune.com', 'books.google.com', 'books.google.com', 'books.google.com', 'taxpaisa.com', 'www.algebra.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.curiouscook.com', 'priyadsouza.com', 'www.cambridge.org', 'whc.unesco.org', 'www.factsaboutindia.org', 'religioustolerance.org', 'sanskritdocuments.org', 'www.jstor.org', 'www.cambridge.org', 'indiatogether.org', 'nrn.org', 'www.pewresearch.org', 'www.bhagavad-gita.org', 'esa.un.org', 'www.lowyinstitute.org', 'southasiaanalysis.org', ['the american journal of human genetics '], ['archaeometry '], ['philosophy east and west '], ['the american journal of human genetics '], ['nature ', 'nature.com '], [' the journal of asian studies'], ['pacific affairs ']]",7564733,Allow all users (no expiry set),80764,22 October 2006,Cop 663 ,2385,14,2006-10-22,2006-10,2006
129,129,Turkic peoples,https://en.wikipedia.org/wiki/Turkic_peoples,261,16,"['10.1017/ehs.2020.11', '10.1017/ehs.2020.4', '10.1016/j.ara.2020.100177', '10.1086/377005', '10.2307/599159', '10.13173/centasiaj.59.1-2.0101', '10.1177/0971945818775373', '10.1093/jis/13.1.75', '10.1038/s41586-018-0094-2', '10.1371/journal.pgen.1005068', '10.1163/25898833-12340008', '10.1163/22105832-00702005', '10.3406/syria.1952.4789', 'abs/10.1177/0971945818775373?journalcode=mhja', '10.1163/22105018-12340089', None, None, None, '12858290', None, None, None, None, '29743675', '25898006', None, None, None, None, None, None, None, None, '1180365', None, None, None, None, None, '4405460', None, None, None, None, None]","[['evolutionary human sciences ', '[[cambridge university press'], ['evolutionary human sciences ', '[[cambridge university press'], ['archaeological research in asia ', '[[elsevier'], [' american journal of human genetics '], ['journal of the american oriental society'], ['central asiatic journal'], ['  the medieval history journal '], ['journal of islamic studies ', '[[oxford centre for islamic studies'], ['[[nature ', '[[nature research'], ['[[plos one', '[[plos'], [' international journal of eurasian linguistics'], ['language dynamics and change ', '[[brill publishers'], ['syria '], ['sage '], ['inner asia ', '[[brill publishers']]",18,20,0,65,0,0,142,0.06896551724137931,0.07662835249042145,0.24904214559386972,0.06130268199233716,0.0,0.20689655172413793,15,"['www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.scwra.gov', 'www.cia.gov', 'www.stat.gov', 'byegm.gov', 'www.loc.gov', 'statistica.gov', 'www.cia.gov', 'www.cia.gov', '2001.ukrcensus.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'books.google.com', 'books.google.com', 'books.google.com', 'geocities.com', 'books.google.com', 'books.google.com', 'www.xjass.com', 'books.google.com', 'www.britannica.com', 'education.yahoo.com', 'global.oup.com', 'www.karakalpak.com', 'books.google.com', 'books.google.com', 'www.xjass.com', 'www.britannica.com', 'books.google.com', 'search.eb.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'bartleby.com', 'www.yeniturkiye.com', 'wanfangdata.com', 'books.google.com', 'www.silk-road.com', 'books.google.com', 'www.allaboutturkey.com', 'books.google.com', 'www.britannica.com', 'm.stlamerican.com', 'www.kamat.com', 'english.al-akhbar.com', 'www.eurasianhistory.com', 'books.google.com', 'www.worldatlas.com', 'www.iranica.com', 'www.britannica.com', 'books.google.com', 'www.al-monitor.com', 'books.google.com', 'www.nisanyansozluk.com', 'www.geocities.com', 'books.google.com', 'www.trtworld.com', 'www.geocities.com', 'www.todayszaman.com', 'books.google.com', 'www.xjass.com', 'www.xjass.com', 'www.kroraina.com', 'www.britannica.com', 'books.google.com', 'www.ethnologue.com', 'books.google.com', 'syrianobserver.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'iranica.com', 'www.britannica.com', 'books.google.com', 'minorityrights.org', 'turksoy.org', 'zh.wikisource.org', 'www.rferl.org', 'zh.wikisource.org', 'zh.wikisource.org', 'turksoy.org', 'www.iranicaonline.org', 'www.rferl.org', 'hk.plm.org', 'zh.wikisource.org', 'www.iranicaonline.org', 'zh.wikisource.org', 'ctext.org', 'www.devplan.org', 'www.iranicaonline.org', 'www.iranicaonline.org', 'www.pbs.org', ['evolutionary human sciences ', '[[cambridge university press'], ['evolutionary human sciences ', '[[cambridge university press'], ['archaeological research in asia ', '[[elsevier'], [' american journal of human genetics '], ['journal of the american oriental society'], ['central asiatic journal'], ['  the medieval history journal '], ['journal of islamic studies ', '[[oxford centre for islamic studies'], ['[[nature ', '[[nature research'], ['[[plos one', '[[plos'], [' international journal of eurasian linguistics'], ['language dynamics and change ', '[[brill publishers'], ['syria '], ['sage '], ['inner asia ', '[[brill publishers']]",44740,Require autoconfirmed or confirmed access (no expiry set),159793,9 November 2001,H. Jonat~enwiki ,5502,25,2001-11-09,2001-11,2001
130,130,Yoruba people,https://en.wikipedia.org/wiki/Yoruba_people,271,24,"['10.1525/ae.1977.4.4.02a00020', '10.1016/j.ajhg.2020.10.010', '10.1038/ncomms7596', '10.1093/acrefore/9780190277734.013.371', '10.1375/1369052023009', '10.1080/0015587x.1959.9717164', '10.1111/j.1471-0528.1960.tb09255.x', '10.1017/s0021853700004035', '10.1057/9781137486431.0006', '10.1007/978-94-6300-121-2_7', '10.1515/9783110860924-008', '10.4314/afrrev.v4i3.60187', '10.4314/afrrev.v3i2.43614', '10.1017/upo9781580466622.002', '10.1017/s0021853700009312', '10.1017/cbo9781107286252.011', '10.20534/eja-16-1-36-45', '10.1017/s0001972017000900', '10.14207/ejsd.2016.v5n1p63', '10.1086/203234', '10.1080/0972639x.2004.11886508', '10.1093/afraf/adw035', '10.1038/nature13997', '10.1126/science.aay5012', None, '33321100', '25803618', None, '11931691', None, '13757217', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, '25470054', '32193295', None, '7820629', '4374169', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, '4297536', '7115999']","[['american ethnologist'], [' ajhg '], ['nature communications '], ['oxford university press'], ['twin research '], ['folklore '], ['bjog'], ['the journal of african history '], ['palgrave macmillan'], ['sensepublishers'], ['de gruyter'], ['african research review'], ['african research review '], ['boydell and brewer limited'], ['journal of african history'], ['cambridge university press'], ['european journal of arts'], ['africa '], ['european journal of sustainable development'], ['current anthropology '], ['studies of tribes and tribals'], ['african affairs '], ['[[nature '], ['science']]",20,4,0,150,0,0,74,0.07380073800738007,0.014760147601476014,0.5535055350553506,0.08856088560885608,0.0,0.17712177121771217,24,"['files.eric.ed.gov', 'data.census.gov', 'www.nps.gov', 'www.cia.gov', 'omojuwa.com', 'books.google.com', 'books.google.com', 'books.google.com', 'raceandhistory.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.google.com', 'books.google.com', 'www.google.com', 'www.google.com', 'beegeagle.wordpress.com', 'www.google.com', 'www.flickr.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'www.coastalnews.com', 'books.google.com', 'books.google.com', 'www.premiumtimesng.com', 'books.google.com', 'www.pmnewsnigeria.com', 'www.google.com', 'www.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'nigeriaworld.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.google.com', 'books.google.com', 'www.ralaran.com', 'www.google.com', 'books.google.com', 'www.google.com', 'grin.com', 'www.jolome.com', 'www.noorimages.com', 'www.mynewswatchtimesng.com', 'www.google.com', 'www.lagbaja.com', 'lulu.com', 'www.google.com', 'books.google.com', 'www.jolome.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.google.com', 'britannica.com', 'books.google.com', 'books.google.com', 'www.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.google.com', 'www.google.com', 'books.google.com', 'books.google.com', 'allafrica.com', 'www.spyghana.com', 'blogdesproductions.wordpress.com', 'books.google.com', 'www.scribd.com', 'books.google.com', 'www.google.com', 'encarta.msn.com', 'books.google.com', 'books.google.com', 'books.google.com', 'academic.oup.com', 'www.google.com', 'www.google.com', 'books.google.com', 'books.google.com', 'www.google.com', 'books.google.com', 'www.cnn.com', 'books.google.com', 'www.post-gazette.com', 'www.jpanafrican.com', 'artsandculture.google.com', 'www.google.com', 'www.imodara.com', 'www.graphic.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.google.com', 'books.google.com', 'www.bbc.com', 'nairametrics.com', 'www.google.com', 'www.google.com', 'books.google.com', 'www.google.com', 'www.aboutlagos.com', 'fashion-history.lovetoknow.com', 'punchng.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.kingdomsofnigeria.com', 'books.google.com', 'rateyourmusic.com', 'books.google.com', 'books.google.com', 'www.imodara.com', 'www.jolome.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.urpress.com', 'books.google.com', 'books.google.com', 'yorupedia.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'nigerianfinder.com', 'www.descarga.com', 'allafrica.com', 'tribuneonlineng.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'unpo.org', 'www.templeoduduwa.org', 'www.yorubaalliance.org', 'escholarship.org', 'unpo.org', 'www.wdl.org', 'www.sciencemag.org', 'www.metmuseum.org', 'international.ipums.org', 'www.jstor.org', 'www.jstor.org', 'www.revistatopoi.org', 'eleda.org', 'www.ekimogundescendant.org', 'www.peoplegroups.org', 'access.thebrightcontinent.org', 'www.fao.org', 'www.peoplegroups.org', 'www.jstor.org', 'globalsecurity.org', ['american ethnologist'], [' ajhg '], ['nature communications '], ['oxford university press'], ['twin research '], ['folklore '], ['bjog'], ['the journal of african history '], ['palgrave macmillan'], ['sensepublishers'], ['de gruyter'], ['african research review'], ['african research review '], ['boydell and brewer limited'], ['journal of african history'], ['cambridge university press'], ['european journal of arts'], ['africa '], ['european journal of sustainable development'], ['current anthropology '], ['studies of tribes and tribals'], ['african affairs '], ['[[nature '], ['science']]",19996678,Allow all users (no expiry set),164206,23 October 2001,130.60.139.xxx ,5404,29,2001-10-23,2001-10,2001
131,131,Zimbabwe,https://en.wikipedia.org/wiki/Zimbabwe,357,13,"['10.1016/s0277-9536(99)00110-0', '10.1038/s41467-020-19493-3', '10.2307/3336358', '10.2307/3889033', '10.2307/219092', '10.1016/s0305-750x(97)00019-3', '10.1016/s0167-8809(99)00156-5', '10.1080/0163660x.2021.1934997', '10.15700/saje.v29n2a259', '10.1093/biosci/bix014', '10.1353/hrq.2010.0030', '10.4102/ve.v36i2.1438', '10.1080/136023699373774', '10414831', '33293507', None, None, None, None, None, None, None, '28608869', None, None, None, None, '7723057', None, None, None, None, None, None, None, '5451287', None, None, None]","[['soc. sci. med.'], ['nature communications'], ['african arts'], ['the south african archaeological bulletin'], ['the international journal of african historical studies'], ['world development'], ['agriculture'], ['the washington quarterly'], ['south african journal of education'], ['bioscience'], ['human rights quarterly'], ['verbum et ecclesia'], [' journal of architecture']]",82,14,0,110,0,6,135,0.22969187675070027,0.0392156862745098,0.3081232492997199,0.036414565826330535,0.0,0.30532212885154064,13,"['www.mod.gov', 'www.parlzim.gov', 'www.mod.gov', 'www.gov', '2001-2009.state.gov', 'www.gov', 'www.gov', 'www.parlzim.gov', 'www.parlzim.gov', 'www.cia.gov', 'www.parlzim.gov', 'harare.usembassy.gov', '2009-2017.state.gov', '2001-2009.state.gov', 'news.google.com', 'www.everycrsreport.com', 'wwp.greenwichmeantime.com', 'www.upi.com', 'www.bloomberg.com', 'www.britannica.com', 'msnbc.com', 'www.africanews.com', 'www.superxv.com', 'www.reuters.com', 'theafricaneconomist.com', 'www.nytimes.com', 'newsofhesouth.com', 'www.infoplease.com', 'www.reuters.com', 'www.cnn.com', 'encarta.msn.com', 'www.reuters.com', 'www.hrforumzim.com', 'www.highbeam.com', 'www.kitco.com', 'www.hrforumzim.com', 'edition.cnn.com', 'www.reuters.com', 'smattgeeksmedia.com', 'www.europeansanctions.com', 'www.sabcnews.com', 'psmag.com', 'ir.imarainvestor.com', 'www.zimbabwedefence.com', 'africareview.com', 'www.dw.com', 'archives.cnn.com', 'books.google.com', 'www.pressreference.com', 'www.sabcnews.com', 'www.newzimbabwe.com', 'allafrica.com', 'www.reuters.com', 'www.zimbabwedefence.com', 'zimbabwemetro.com', 'biztechafrica.com', 'edition.cnn.com', 'www.google.com', 'www.newsdeeply.com', 'www.bbc.com', 'www.cnn.com', 'www.nytimes.com', 'about.com', 'www.cnn.com', 'zimbabwe-today.com', 'af.reuters.com', 'allafrica.com', 'www.reuters.com', 'www.aljazeera.com', 'www.nybooks.com', 'zambuko.com', 'sportsillustrated.cnn.com', 'www.bbc.com', 'www.sokwanele.com', 'af.reuters.com', 'www.newzimbabwe.com', 'ed.ted.com', 'www.reuters.com', 'www.somalipress.com', 'www.historytoday.com', 'africa.reuters.com', 'www.economist.com', 'query.nytimes.com', 'infoplease.com', 'news.sky.com', 'www.burnhamkingofscouts.com', 'www.cnn.com', 'richardknight.homestead.com', 'africantears.netfirms.com', 'gapadventures.com', 'www.voazimbabwe.com', 'www.washingtonpost.com', 'zimbabwejournalists.com', 'www.csmonitor.com', 'karaart.com', 'www.britannica.com', 'www.time.com', 'www.reuters.com', 'news.nationalgeographic.com', 'www.talkzimbabwe.com', 'www.reuters.com', 'www.peakbagger.com', 'zimbabwemetro.com', 'www.gapadventures.com', 'archives.cnn.com', 'money.cnn.com', 'www.britannica.com', 'www.voanews.com', 'www.thezimbabwemail.com', 'www.economist.com', 'zwnews.com', 'www.trtworld.com', 'books.google.com', 'www.newzimbabwe.com', 'www.smh.com', 'www.usatoday.com', 'www.thesculpturepark.com', 'www.sabcnews.com', 'www.cnn.com', 'www.washingtonpost.com', 'www.foxnews.com', 'members.fortunecity.com', 'www.britannica.com', 'biztechafrica.com', 'www.sahistory.org', 'rsf.org', 'www.wttc.org', 'www.eisa.org', 'cpj.org', 'data.worldbank.org', 'www.radionetherlandsarchives.org', 'www.ifex.org', 'www.undp.org', 'www.eisa.org', 'www.internal-displacement.org', 'www.worldbank.org', 'web.amnesty.org', 'www.cato.org', 'www.zw.one.un.org', 'africanarguments.org', 'www.unhcr.org', 'thecommonwealth.org', 'www.icrisat.org', 'www.hrw.org', 'unesdoc.unesco.org', 'hrw.org', 'www.pewforum.org', 'www.sahistory.org', 'eiard.org', 'www.cgdev.org', 'www.zw.one.un.org', 'www.icrc.org', 'news.un.org', 'www.hrw.org', 'unesdoc.unesco.org', 'www.eisa.org', 'www.undp.org', 'www.undp.org', 'www.irinnews.org', 'npr.org', 'zimbabwe.poetryinternationalweb.org', 'www.sahistory.org', 'www.unocha.org', 'countrystat.org', 'www.mantleplumes.org', 'www.unfpa.org', 'irinnews.org', 'www.humanrightsfirst.org', 'worldrugby.org', 'www.unocha.org', 'www.fina.org', 'adventistatlas.org', 'media.ifrc.org', 'www.sahistory.org', 'esa.un.org', 'www.hrw.org', 'www.radionetherlandsarchives.org', 'www.un.org', 'www.undp.org', 'www.fina.org', 'www.nrzam.org', 'www.chathamhouse.org', 'www.avert.org', 'www.harare.unesco.org', 'www.unaids.org', 'unstats.un.org', 'www.hrw.org', 'news.amnesty.org', 'www.fao.org', 'www.unaids.org', 'www.imf.org', 'freedomhouse.org', 'issafrica.org', 'www.zw.one.un.org', 'www.zw.one.un.org', 'hdr.undp.org', 'victoriafallstourism.org', 'heritage.org', 'www.undp.org', 'zimeye.org', 'wsp.org', 'ilga.org', 'www.fao.org', 'www.undp.org', 'www.jstor.org', 'zimbabwe.unfpa.org', ['soc. sci. med.'], ['nature communications'], ['african arts'], ['the south african archaeological bulletin'], ['the international journal of african historical studies'], ['world development'], ['agriculture'], ['the washington quarterly'], ['south african journal of education'], ['bioscience'], ['human rights quarterly'], ['verbum et ecclesia'], [' journal of architecture']]",34399,Require administrator access (no expiry set),225234,13 March 2001,JimboWales ,12220,38,2001-03-13,2001-03,2001
132,132,Venice,https://en.wikipedia.org/wiki/Venice,197,3,"['10.1111/j.1477-4658.1999.tb00064.x', '10.1017/aaq.2021.38', '10.1484/j.viator.2.301504', None, None, None, None, None, None]","[['renaissance studies ', '[[wiley '], ['american antiquity '], ['viator ']]",20,1,0,73,0,8,92,0.10152284263959391,0.005076142131979695,0.37055837563451777,0.015228426395939087,0.0,0.1218274111675127,3,"['www.mit.gov', 'www.huffingtonpost.com', 'britannica.com', 'time.com', 'books.google.com', 'www.sci-news.com', 'www.forbes.com', 'www.moovitapp.com', 'www.smithsonianmag.com', 'news.sky.com', 'bbc.com', 'www.studyabroad.com', 'www.ibtimes.com', 'live.com', 'www.bbc.com', 'arthistory.about.com', 'www.moovitapp.com', 'www.bbc.com', 'www.ft.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.bbc.com', 'www.cnn.com', 'www.nytimes.com', 'www.latimes.com', 'www.theverge.com', 'www.reuters.com', 'www.cnn.com', 'veneziaautentica.com', 'books.google.com', 'www.nytimes.com', 'livescience.com', 'www.ricksteves.com', 'www.com', 'dstandish.com', 'books.google.com', 'veneziaautentica.com', 'money.cnn.com', 'www.com', 'news.artnet.com', 'www.ilsole24ore.com', 'time.com', 'www.hotelsantelena.com', 'www.etymonline.com', 'www.washingtonpost.com', 'news.nationalgeographic.com', 'books.google.com', 'books.google.com', 'www.cruisetradenews.com', 'www.ikonlondonmagazine.com', 'www.britannica.com', 'www.nytimes.com', 'www.com', 'www.lonelyplanet.com', 'www.themeshnews.com', 'worldchacha.com', 'live.com', 'www.washingtonpost.com', 'www.weather-atlas.com', 'www.newsweek.com', 'www.nytimes.com', 'www.euronews.com', 'www.reuters.com', 'www.forbes.com', 'europeforvisitors.com', 'edition.cnn.com', 'www.cruisearabiaonline.com', 'britannica.com', 'venicegondola.com', 'www.anglenews.com', 'www.hollywoodreporter.com', 'books.google.com', 'books.google.com', 'www.nationalgallery.org', 'webexhibits.org', 'www.seatemperature.org', 'catholic-hierarchy.org', 'labiennale.org', 'www.npr.org', 'labiennale.org', 'weareherevenice.org', 'www.treesforlife.org', 'aboutvenice.org', 'whc.unesco.org', 'www.pbs.org', 'npr.org', 'dbs.bh.org', 'iranicaonline.org', 'www.jewishvirtuallibrary.org', 'www.cvni.org', 'www.seatemperature.org', 'www.univiu.org', 'www.pbs.org', ['renaissance studies ', '[[wiley '], ['american antiquity '], ['viator ']]",32616,Require administrator access (no expiry set),164028,6 October 2001,Trimalchio ,9353,14,2001-10-06,2001-10,2001
133,133,Turkey,https://en.wikipedia.org/wiki/Turkey,545,15,"['10.1016/j.geothermics.2005.09.003', '10.1016/j.apr.2020.08.011', '10.2307/632236', '10.1017/npt.2018.7', '10.1017/s0020743800063819', '10.1126/science.303.5662.1323', '10.1080/00905990500504871', '10.18452/3090', '10.1007/978-3-030-03515-0_36', '10.2307/3258667', '10.1093/hgs/12.3.393', '10.1080/01419870701491937', '10.1080/13537110208428662', '10.1080/14623520801950820', None, None, None, None, None, '14988549', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None]","[['geothermics'], ['atmospheric pollution research'], ['the journal of hellenic studies'], ['new perspectives on turkey'], ['international journal of middle east studies '], ['science'], ['[[nationalities papers'], ['humboldt-universität zu berlin'], ['springer international publishing'], ['the metropolitan museum of art bulletin'], ['holocaust and genocide studies'], ['ethnic and racial studies'], ['nationalism and ethnic politics', 'yale university'], ['journal of genocide research']]",86,61,0,192,0,6,186,0.1577981651376147,0.11192660550458716,0.3522935779816514,0.027522935779816515,0.0,0.29724770642201837,14,"['www.cia.gov', 'www.mfa.gov', 'mfa.gov', 'www.yok.gov', 'www.resmigazete.gov', 'tubitak.gov', 'www.resmigazete.gov', 'www.mfa.gov', 'www.cia.gov', 'www.anayasa.gov', 'envanter.gov', 'www.turkiyeburslari.gov', 'www.taek.gov', 'www.dmi.gov', 'www.tccb.gov', 'www.state.gov', 'kvmgm.ktb.gov', 'www.cia.gov', 'mfa.gov', 'www.turkstat.gov', 'data.tuik.gov', 'www.kultur.gov', 'www.tbmm.gov', 'www.dhmi.gov', 'www.e-icisleri.gov', 'www.rtuk.gov', 'www.mfa.gov', 'mfa.gov', 'mfa.gov', 'data.tuik.gov', 'www.abgs.gov', 'mfa.gov', 'mfa.gov', 'www.studyinturkey.gov', 'www.kgm.gov', 'state.gov', 'uhdigm.adalet.gov', 'www.kultur.gov', 'lcweb2.loc.gov', 'tuba.gov', 'cia.gov', 'www.ssm.gov', 'www.anayasa.gov', 'milliparklar.gov', 'lcweb2.loc.gov', 'tcmb.gov', 'mfa.gov', 'www.mfa.gov', 'mfa.gov', 'global.tbmm.gov', 'www.cia.gov', 'www.ysk.gov', 'www.ab.gov', 'mfa.gov', 'www.anayasa.gov', 'yigm.kulturturizm.gov', 'www.anayasa.gov', 'hizlitren.tcdd.gov', 'www.turkstat.gov', 'www.die.gov', 'justice.gov', 'books.google.com', 'www.worldatlas.com', 'edition.cnn.com', 'www.aa.com', 'www.hurriyetdailynews.com', 'kirkpinar.com', 'milliyet.com', 'bbc.com', 'www.ethnologue.com', 'www.dw.com', 'www.bloomberg.com', 'www.konda.com', 'worldhistory.byethost8.com', 'www.dw.com', 'www.trtworld.com', 'www.bbc.com', 'aljazeera.com', 'allaboutturkey.com', 'books.google.com', 'hurarsiv.hurriyet.com', 'hurriyetdailynews.com', 'www.bloomberg.com', 'gazeteciler.com', 'aa.com', 'www.climatechangenews.com', 'latitude.blogs.nytimes.com', 'books.google.com', 'www.hurriyetdailynews.com', 'www.gercekgundem.com', 'books.google.com', 'www.bbc.com', 'books.google.com', 'www.ebrd.com', 'books.google.com', 'www.hurriyet.com', 'www.ft.com', 'books.google.com', 'www.al-monitor.com', 'tarkandeluxe.blogspot.com', 'global.britannica.com', 'www.gazeteduvar.com', 'igairport.com', 'books.google.com', 'www.reuters.com', 'www.newsweek.com', 'assets.new.siemens.com', 'jewishencyclopedia.com', 'allaboutturkey.com', 'books.google.com', 'www.sozcu.com', 'foodbycountry.com', 'www.sacred-texts.com', 'www.oxfordreference.com', 'books.google.com', 'www.britannica.com', 't24.com', 'thedefensepost.com', 'www.bbc.com', 'www.dailysabah.com', 'books.google.com', 'books.google.com', 'www.ibtimes.com', 'www.bbc.com', 'digiday.com', 'www.trtworld.com', 'turkresmi.com', 'www.ipsosglobaltrends.com', 'www.dw.com', 'emreozgur.com', 'www.reuters.com', 'ancienthistory.about.com', 'www.ncturkishfestival.com', 'www.dailysabah.com', 'www.reuters.com', 'books.google.com', 'www.economist.com', 'www.ntv.com', 'books.google.com', 'books.google.com', 'www.karalahana.com', 'english.peopledaily.com', 'europe.newsweek.com', 'bloomberg.com', 'www.nytimes.com', 'www.bbc.com', 'www.reuters.com', 'www.reuters.com', 'fibaeurope.com', 'books.google.com', 'www.aa.com', 'www.psychiatrictimes.com', 'www.saudiaramcoworld.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.defensenews.com', 'dolmabahcepalace.com', 'atelyemim.com', 'www.hurriyet.com', 'www.hurriyetdailynews.com', 'www.trthaber.com', 'www.hurriyetdailynews.com', 'aksiyon.com', 'www.bloomsbury.com', 'books.google.com', 'books.google.com', 'www.dailysabah.com', 'biblehub.com', 'www.nytimes.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'www.businessweek.com', 'www.sozcu.com', 'www.nytimes.com', 'www.topuniversities.com', 'investor.turkishairlines.com', 'www.aa.com', 'www.springer.com', 'www.hurriyet.com', 'books.google.com', 'turkeyscholarship.com', 'books.google.com', 'www.defensenews.com', 'akkunpp.com', 'ahvalnews.com', 'go.euromonitor.com', 'arsiv.ntvmsnbc.com', 'books.google.com', 'www.reuters.com', 'www.iphs2010.com', 'www.reuters.com', 'books.google.com', 'books.google.com', 'www.al-monitor.com', 'www.dw.com', 'simitcay.com', 'www.aljazeera.com', 'www.hurriyetdailynews.com', 'www.msn.com', 'uefa.com', 'cadde.milliyet.com', 'fibaeurope.com', 'britannica.com', 'britannica.com', 'www.lesartsturcs.com', 'www.goturkey.com', 'blog.oup.com', 'books.google.com', 'www.reuters.com', 'www.bbc.com', 'www.reuters.com', 'www.cnn.com', 'www.reuters.com', 'www.dailysabah.com', 'www.dailysabah.com', 'foreignpolicy.com', 'www.hurriyetdailynews.com', 'www.hurriyetdailynews.com', 'www.trtworld.com', 'britannica.com', 'turkeypurge.com', 'bloomberg.com', 'www.nytimes.com', 'books.google.com', 'www.newsweek.com', 'global.britannica.com', 'www.al-monitor.com', 'www.aljazeera.com', 'www.nytimes.com', 'dw.com', 'books.google.com', 'books.google.com', 'www.al-monitor.com', 'www.dailysabah.com', 'www.reuters.com', 'edition.cnn.com', 'www.trtworld.com', 'gateofturkey.com', 'www.euronews.com', 'allaboutturkey.com', 'books.google.com', 'books.google.com', 'www.dw.com', 'www.cnbc.com', 'www.ipsos-na.com', 'www.foreignaffairs.com', 'www.reuters.com', 'www.washingtonpost.com', 'books.google.com', 'hurriyet.com', 'books.google.com', 'freedomhouse.org', 'www.turkishculture.org', 'fas.org', 'esn.org', 'mimarlikmuzesi.org', 'hdr.undp.org', 'en.efesbasket.org', 'islamansiklopedisi.org', 'data2.unhcr.org', 'cpj.org', 'tvf.org', 'www.nrdc.org', 'archmuseum.org', 'data.worldbank.org', 'www-wds.worldbank.org', 'www.turks.org', 'www.worldhistory.org', 'www.transparency.org', 'stats.oecd.org', 'data.worldbank.org', 'www.shura.org', 'www.iranicaonline.org', 'freemuse.org', 'catholic-hierarchy.org', 'www.worldhistory.org', 'esiweb.org', 'turkishculture.org', 'christiancentury.org', 'bianet.org', 'whc.unesco.org', 'esa.un.org', 'www.turkishculture.org', 'tff.org', 'iucn.org', 'www.imf.org', 'cpj.org', 'fenerbahce.org', 'bianet.org', 'unhcr.org', 'www.bianet.org', 'www.uncyprustalks.org', 'cpj.org', 'www.wes.org', 'carbontracker.org', 'www-wds.worldbank.org', 'www.worldhistory.org', 'www.worldbank.org', 'eczacibasisporkulubu.org', 'www.oecd.org', 'unstats.un.org', 'www.meforum.org', 'www.studyinturkey.org', 'refworld.org', 'www.khrp.org', 'www.iea.org', 'wayback.archive-it.org', 'www.unesco.org', 'www.jewishdatabank.org', 'www.jewishvirtuallibrary.org', 'www.americansephardifederation.org', 'archnet.org', 'www.unhcr.org', 'newsroom.churchofjesuschrist.org', 'www.shura.org', 'www.aina.org', 'turkishculture.org', 'peter.mackenzie.org', 'www.archaeology.org', 'www.metmuseum.org', 'www.minorityrights.org', 'www.pewforum.org', 'ancienthistorybulletin.org', 'tesev.org', 'data.worldbank.org', 'www.oecd.org', 'en.efesbasket.org', 'www.carnegieendowment.org', 'en.wikipedia.org', 'www.shura.org', 'www.metmuseum.org', 'www.un.org', 'pulitzercenter.org', 'turkishculture.org', 'weekly.ahram.org', 'globalheritagefund.org', 'www.unesco.org', ['geothermics'], ['atmospheric pollution research'], ['the journal of hellenic studies'], ['new perspectives on turkey'], ['international journal of middle east studies '], ['science'], ['[[nationalities papers'], ['humboldt-universität zu berlin'], ['springer international publishing'], ['the metropolitan museum of art bulletin'], ['holocaust and genocide studies'], ['ethnic and racial studies'], ['nationalism and ethnic politics', 'yale university'], ['journal of genocide research']]",11125639,Require administrator access (no expiry set),299951,2 September 2001,Zundark ,21996,32,2001-09-02,2001-09,2001
134,134,Rajasthani people,https://en.wikipedia.org/wiki/Rajasthani_people,62,1,"['10.24321/2456.0510.201808', None, None]",[['anusanadhan']],0,1,0,17,0,0,43,0.0,0.016129032258064516,0.27419354838709675,0.016129032258064516,0.0,0.03225806451612903,1,"['www.rajasthan.gov', 'www.britannica.com', 'www.google.com', 'www.bharatonline.com', 'm.timesofindia.com', 'books.google.com', 'books.google.com', 'books.google.com', 'journeymart.com', 'economictimes.indiatimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'travel-in-rajasthan.com', 'travel-in-rajasthan.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', ['anusanadhan']]",23041891,Allow all users (no expiry set),39646,1 June 2009,Saimdusan ,1019,32,2009-06-01,2009-06,2009
135,135,Fricassee,https://en.wikipedia.org/wiki/Fricassee,19,0,[],[],0,0,0,8,0,0,11,0.0,0.0,0.42105263157894735,0.0,0.0,0.0,0,"['www.etymonline.com', 'www.lexico.com', 'www.lafayettetravel.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.elboricua.com']",9125820,Allow all users (no expiry set),9607,26 January 2007,Bigtrick ,232,5,2007-01-26,2007-01,2007
136,136,Uttar Pradesh,https://en.wikipedia.org/wiki/Uttar_Pradesh,303,4,"['10.4103/0019-557x.138624', '10.1017/s0026749x00015092', '10.1007/bf02704749', '10.1016/j.quascirev.2007.11.001', '25116823', None, '11779962', None, None, None, None, None]","[['indian journal of public health '], ['modern asian studies'], ['journal of biosciences ', '[[indian academy of sciences'], ['quaternary science reviews']]",21,55,0,140,0,0,83,0.06930693069306931,0.18151815181518152,0.46204620462046203,0.013201320132013201,0.0,0.264026402640264,4,"['www.censusindia.gov', 'www.uptourism.gov', 'uphome.gov', 'upforest.gov', 'amrut.gov', 'www.imd.gov', 'ncrb.gov', 'censusindia.gov', 'www.upgovernor.gov', 'www.imd.gov', 'censusindia.gov', 'upforest.gov', 'uptourism.gov', 'www.up.gov', 'uppolice.gov', 'www.imd.gov', 'up.gov', 'amrut.gov', 'www.uptourism.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'www.niti.gov', 'www.ner.indianrailways.gov', 'www.imd.gov', 'www.archive.india.gov', 'censusmp.gov', 'archive.india.gov', 'upforest.gov', 'upforest.gov', 'censusindia.gov', 'www.farmech.dac.gov', 'www.imd.gov', 'censusindia.gov', 'ncl.gov', 'up.gov', 'censusindia.gov', 'www.trai.gov', 'censusindia.gov', 'pib.gov', 'www.indianrailways.gov', 'www.censusindia.gov', 'idup.gov', 'zsi.gov', 'censusindia.gov', 'ncr.indianrailways.gov', 'www.censusindia.gov', 'up.gov', 'planningcommission.gov', 'niti.gov', 'uplegisassembly.gov', 'www.imd.gov', 'india.gov', 'www.imd.gov', 'uplegisassembly.gov', 'lko.railnet.gov', 'books.google.com', 'timesofindia.indiatimes.com', 'articles.timesofindia.indiatimes.com', 'zeenews.india.com', 'thehaider.com', 'www.up-tourism.com', 'books.google.com', 'www.tehelka.com', 'books.google.com', 'post.jagran.com', 'www.thehindubusinessline.com', 'books.google.com', 'www.firstpost.com', 'www.up-tourism.com', 'economictimes.indiatimes.com', 'www.hindustantimes.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.weather.com', 'books.google.com', 'articles.timesofindia.indiatimes.com', 'www.up-tourism.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'indiansugar.com', 'www.jagranjosh.com', 'paper.hindustantimes.com', 'www.masterplansindia.com', 'rediff.com', 'www.whatisindia.com', 'www.indfy.com', 'zeenews.india.com', 'rediff.com', 'www.hindu.com', 'books.google.com', 'www.greaternoida.com', 'books.google.com', 'www.thesundayindian.com', 'books.google.com', 'fmstations.bharatiyamobile.com', 'economictimes.indiatimes.com', 'economictimes.indiatimes.com', 'economictimes.indiatimes.com', 'www.hindustantimes.com', 'books.google.com', 'books.google.com', 'www.youtube.com', 'in.news.yahoo.com', 'www.hindustantimes.com', 'books.google.com', 'articles.timesofindia.indiatimes.com', 'books.google.com', 'articles.economictimes.indiatimes.com', 'www.hindu.com', 'amsglossary.allenpress.com', 'books.google.com', 'www.thehindubusinessline.com', 'www.newindianexpress.com', 'zeenews.india.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.stick2hockey.com', 'newkerala.com', 'www.ndtv.com', 'economictimes.indiatimes.com', 'www.indiatimes.com', 'www.india-cellular.com', 'www.upfcindia.com', 'www.indianexpress.com', 'www.business-standard.com', 'books.google.com', 'articles.timesofindia.indiatimes.com', 'www.jaypeesports.com', 'www.business-standard.com', 'www.business-standard.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.ethnologue.com', 'www.educationinfoindia.com', 'www.hindustantimes.com', 'www.thehindu.com', 'books.google.com', 'www.hindustantimes.com', 'books.google.com', 'www.upfcindia.com', 'www.hindustantimes.com', 'www.noidaauthorityonline.com', 'books.google.com', 'www.jagranjosh.com', 'www.moneycontrol.com', 'www.ndtv.com', 'www.lexuniverse.com', 'www.jagranjosh.com', 'articles.timesofindia.indiatimes.com', 'www.benaresmusicacademy.com', 'rediff.com', 'www.livemint.com', 'books.google.com', 'books.google.com', 'qz.com', 'www.indianexpress.com', 'books.google.com', 'www.livemint.com', 'sites.google.com', 'www.newindianexpress.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'www.indianexpress.com', 'books.google.com', 'articles.timesofindia.indiatimes.com', 'www.hindustaniclassical.com', 'www.webindia123.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.jagranjosh.com', 'economictimes.indiatimes.com', 'ibnlive.in.com', 'zeenews.india.com', 'articles.timesofindia.indiatimes.com', 'books.google.com', 'www.aljazeera.com', 'www.hindustantimes.com', 'www.mapsofindia.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.deccanherald.com', 'books.google.com', 'news.webindia123.com', 'amsglossary.allenpress.com', 'www.mbauniverse.com', 'books.google.com', 'books.google.com', 'www.hindustantimes.com', 'books.google.com', 'rbidocs.rbi.org', 'www.gecafs.org', 'asci.org', 'www.ibef.org', 'upsbdb.org', 'www.cehat.org', 'www.ibef.org', 'documents.worldbank.org', 'documents.worldbank.org', 'www.janaagraha.org', 'ibef.org', 'ww.orientalbirdclub.org', 'www.worldartswest.org', 'www.prsindia.org', 'www.hindunet.org', 'www.jstor.org', 'www.lawsofindia.org', 'www.fsi.org', 'hdi.globaldatalab.org', 'hdr.undp.org', 'www.rbi.org', ['indian journal of public health '], ['modern asian studies'], ['journal of biosciences ', '[[indian academy of sciences'], ['quaternary science reviews']]",231623,"Require autoconfirmed or confirmed access (18:07, 10 May 2023)",212139,22 May 2003,Caid Raspa ,8211,16,2003-05-22,2003-05,2003
137,137,Russia,https://en.wikipedia.org/wiki/Russia,614,171,"['10.1163/187633106x00186', '10.1017/slr.2018.13', '10.12797/politeja.12.2015.31_2.09', '10.2307/3020237', '10.2307/1174124', '10.2307/898239', '10.1093/musqtl/gdm001', '10.55540/0031-1723.2944', '10.1080/07075332.2009.9641172', '10.1098/rsbm.1977.0004', '10.2307/1836520', '10.1787/d8b068b4-en', '10.1177/0967010602033001006', '10.1093/oxartj/12.1.14', '10.1086/418982', '10.1017/nps.2019.14', '10.2307/3000442', '10.1093/publius/pjl004', '10.5699/slaveasteurorev2.97.2.0227', '10.1038/s41467-020-19493-3', '10.1038/ejhg.2017.117', '10.1093/mq/xiii.1.29', '10.1126/science.aao1807', '10.2307/126593', '10.1086/649363', '10.2307/125254', '10.2307/40202977', '10.1080/00210862.2012.758502', '10.1093/wbro/13.1.37', '10.2307/3049132', '10.1080/09668130500401715', '10.2307/377158', '10.2307/20029588', '10.2307/2137719', '10.2307/129919', '10.1016/j.ygeno.2019.03.007', '10.2307/20030251', '10.2307/j.ctt21h4wkb.15', '10.2139/ssrn.1333553', '10.1177/030631278101100201', '10.7592/fejf2015.62', '10.2307/3679044', '10.2307/127655', '10.1098/rsbm.1936.0001', '10.1038/35006625', '10.1080/14623528.2020.1834741', '10.1179/sic.2009.54.1.12', '10.2307/127159', '10.2307/2320506', '10.1080/01436599714911', '10.2307/204825', '10.1177/002200948702200203', '10.1080/00905992.2014.998043', '10.2307/25587683', '10.1353/not.2002.0113', '10.1017/s0960777309005074', '10.1177/000271623920300106', '10.2307/1347433', '10.1136/jech-2020-213885', '10.1353/jwh.2013.0031', '10.2861/664907', '10.1163/187633186x00016', '10.1093/jdh/10.2.177', '10.1111/j.1540-5893.2008.00333.x', '10.1080/09668139808412522', '10.1038/sdata.2018.214', '10.1080/09668139708412462', '10.2307/125859', '10.1175/1520-0469(1971)028<0263:slovot>2.0.co;2', '10.1038/s41586-018-0870-z', '10.2307/1478046', '10.1525/as.2017.57.1.93', '10.1016/j.postcomstud.2012.12.010', '10.2307/2952082', '10.2307/309128', '10.1080/00085006.2003.11092333', '10.1017/s153759270505005x', '10.1017/cbo9780511524028.002', '10.1353/not.2011.0120', '10.11610/connections.14.2.01', '10.1257/0895330053147949', '10.2307/2534597', '10.1017/s0020818300004859', None, '10.1159/000443331', '10.5129/001041518822704872', '10.1080/00045608.2010.534713', '10.1163/18763324-04602003', '10.18111/wtobarometereng', '10.2307/2708192', '10.1093/alcalc/34.6.824', '10.1016/s0140-6736(19)32265-2', '10.1007/bf00717701', '10.1038/s41566-019-0525-0', '10.2307/990455', '10.1038/nphoton.2007.34', '10.1163/1571811031310738', '10.2307/125154', '10.1177/002200949703200303', '10.2307/965578', '10.1038/35092552', '10.2307/2534584', '10.5038/1944-0472.12.2.1727', '10.1080/07075332.1989.9640530', '10.1093/past/129.1.168', '10.1093/ml/l.1.153', '10.1787/0b8f90e9-en', '10.1080/09668139408412190', '10.2307/1503933', '10.2307/127973', '10.1057/jird.2008.7', '10.1353/nlh.1998.0040', '10.2307/128091', '10.3390/ijerph16101848', '10.1016/j.postcomstud.2015.12.002', '10.2307/27757115', '10.1177/002200948802300207', '10.2307/1945179', '10.1146/annurev-linguist-030514-124812', '10.2307/126692', '10.1080/08911916.2000.11644017', '10.21273/hortsci.50.6.772', '10.1080/0966813052000314101', '10.1137/070702710', '10.1111/j.1743-8594.2006.00023.x', '10.11610/connections.14.4.08', '10.1086/244076', '10.1038/scientificamerican0897-72', '10.1080/00085006.1984.11091776', '10.2307/2644534', '10.1186/s12889-020-08464-4', '10.2307/1835935', '10.1558/jsrnc.39114', '10.2307/2496635', '10.2307/2953371', '10.1017/s0034670500043965', '10.2307/2491790', '10.1051/shsconf/202111005011', '10.2307/20040512', '10.1136/bmj.1.5113.1', '10.2307/2493225', '10.1080/07075332.1994.9640668', '10.1353/jhi.2015.0028', '10.2307/1833615', '10.1080/09668130903506847', '10.2307/2709278', '10.1080/00029890.2009.11920920', '10.1163/15730352-bja10003', '10.1191/0968344503wh260oa', '10.2307/1945868', '10.1080/00085006.1980.11091635', '10.1093/jaarel/lxii.3.747', '10.2307/1844479', '10.1016/j.quaint.2015.10.032', '10.5840/monist192737121', '10.2307/126075', '10.1016/j.jhevol.2018.11.012', '10.2307/125968', '10.1177/0022009403038001961', '10.5840/raven2012197', '10.2307/20433998', '10.1057/pol.2009.18', '10.1016/j.mayocp.2011.11.003', '10.1038/d41586-018-06004-0', '10.3366/e096813610800037x', '10.1038/nature13810', '10.2307/987741', '10.1163/18763316-04301004', '10.1080/01434632.2010.536237', '10.2307/210882', '10.17104/1611-8944-2015-4-458', None, None, None, None, None, None, None, None, None, '11615738', None, None, None, None, None, None, None, None, None, '33293507', '28905876', None, '28982795', None, None, None, None, None, None, None, None, None, None, None, None, '30902755', None, None, None, None, None, None, None, None, '10761915', None, None, None, None, None, None, None, None, None, None, None, None, None, '32414935', None, None, None, None, None, None, '30375988', None, None, None, '30700871', None, None, None, None, None, None, None, None, None, None, None, None, None, None, '26836137', None, None, None, None, None, '10659717', '31591968', None, None, None, None, None, None, None, None, '11544525', None, None, None, None, None, None, '12288331', None, None, None, None, None, '31137705', None, None, '11617302', None, None, None, None, None, None, None, None, None, None, None, None, None, '32293365', None, None, None, None, None, None, None, None, '13608066', None, None, '26522713', None, None, None, None, None, None, None, None, None, None, None, None, None, '30777356', None, None, None, None, None, '22212977', '30135540', None, '25341783', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, '7723057', '5602018', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, '7577103', None, None, None, None, None, None, '6207062', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, '99322', '6738810', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, '6571548', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, '7092419', None, None, None, None, None, None, None, None, '1992347', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, '3498096', None, None, '4753769', None, None, None, None, None]","[['[[russian history '], ['[[cambridge university press', '[[slavic review'], ['politeja ', 'księgarnia akademicka '], ['[[the slavonic and east european review', '[[cambridge university press'], ['proceedings of the academy of political science ', '[[the academy of political science'], ['[[notes ', '[[music library association'], ['[[oxford university press', 'the musical quarterly'], ['[[parameters '], ['[[taylor ', '[[the international history review'], ['[[biographical memoirs of fellows of the royal society'], ['[[the american historical review', '[[oxford university press'], ['[[oecd'], ['[[sage publishing', '[[security dialogue'], ['[[oxford university press', 'oxford art journal'], ['the [[university of chicago press', '[[the quarterly review of biology'], ['[[nationalities papers'], ['[[slavic review', '[[cambridge university press'], ['[[oxford university press', '[[publius '], ['[[the slavonic and east european review', '[[modern humanities research association'], ['nature communications '], ['[[european journal of human genetics'], ['[[oxford university press', '[[the musical quarterly'], ['science '], ['[[the russian review'], ['the [[university of chicago press', '[[osiris'], ['[[the russian review', '[[wiley '], ['[[canadian international council', '[[sage publishing'], ['[[iranian studies', '[[taylor '], ['the world bank research observer ', '[[oxford university press'], ['caa ', '[[the art bulletin'], ['[[europe-asia studies'], ['[[college english', '[[national council of teachers of english'], ['[[council on foreign relations', '[[foreign affairs'], ['[[population and development review', '[[population council'], ['[[the russian review'], ['genomics ', '[[elsevier'], ['[[council on foreign relations', '[[foreign affairs'], ['[[academic studies press'], ['[[centre for european policy studies'], ['[[sage publishing', '[[social studies of science'], ['folklore'], ['[[royal historical society', '[[cambridge university press'], ['[[the russian review'], ['[[royal society', '[[obituary notices of fellows of the royal society'], [' [[nature '], ['[[journal of genocide research'], ['studies in conservation ', '[[taylor '], ['[[the russian review'], ['[[taylor ', '[[the american mathematical monthly'], ['[[third world quarterly', '[[taylor '], ['[[the journal of interdisciplinary history', 'the [[mit press'], ['[[journal of contemporary history', '[[sage publishing'], ['[[nationalities papers', '[[cambridge university press'], ['the art world'], ['[[notes '], ['[[princeton university', '[[contemporary european history'], ['the annals of the [[american academy of political and social science', '[[sage publishing'], ['rocky mountain modern language association ', 'rocky mountain review of language and literature'], ['journal of epidemiology and community health '], ['[[journal of world history', '[[university of hawaiʻi press'], ['[[european parliamentary research service', '[[european parliament'], ['[[russian history ', '[[brill publishers'], ['[[oxford university press', '[[journal of design history'], ['[[law ', '[[wiley '], ['[[taylor ', '[[europe-asia studies'], ['scientific data '], ['[[europe-asia studies', '[[taylor '], ['[[the russian review', '[[wiley '], ['[[academy of sciences of the soviet union', 'journal of the atmospheric sciences'], ['nature '], ['dance studies association ', '[[congress on research in dance'], ['[[university of california press', '[[asian survey'], ['communist and post-communist studies ', '[[university of california press'], ['the american political science review ', '[[american political science association'], [' [[the slavic and east european journal'], ['[[canadian slavonic papers'], ['[[perspectives on politics', '[[american political science association'], ['[[cambridge university press'], ['[[notes ', '[[music library association'], ['connections ', '[[partnership for peace consortium of defense academies and security studies institutes'], ['[[journal of economic perspectives', '[[harvard university'], ['[[brookings papers on economic activity', '[[brookings institution'], ['[[international organization', 'the [[mit press'], ['canadian medical association journal '], ['journal of innate immunity '], ['comparative politics ', '[[city university of new york'], ['[[annals of the association of american geographers', '[[taylor '], ['the soviet and post-soviet review', 'brill'], ['unwto world tourism barometer english version ', '[[world tourism organization'], ['[[university of pennsylvania press', '[[journal of the history of ideas'], ['alcohol and alcoholism '], ['[[the lancet'], ['geojournal '], ['[[nature photonics'], ['[[university of california press', '[[journal of the society of architectural historians'], ['[[nature photonics'], ['international journal on minority and group rights ', '[[brill publishers'], ['[[wiley ', '[[the russian review'], ['[[journal of contemporary history', '[[sage publishing'], ['[[the musical times'], ['nature '], ['[[brookings papers on economic activity'], ['[[journal of strategic security', '[[university of south florida'], ['[[the international history review'], ['[[past ', '[[oxford university press'], ['[[oxford university press', '[[music '], ['[[oecd'], ['[[europe-asia studies'], ['the journal of decorative and propaganda arts ', '[[florida international university'], ['[[the russian review', '[[wiley '], ['journal of international relations and development'], ['[[the johns hopkins university press', ' [[new literary history'], ['[[the russian review', '[[wiley '], ['[[international journal of environmental research and public health'], ['communist and post-communist studies', '[[university of california press'], ['[[university of california press', '[[chymia'], ['[[journal of contemporary history', '[[sage publishing'], ['[[the american political science review', '[[american political science association'], ['annual review of linguistics '], ['[[wiley ', '[[the russian review'], ['[[taylor ', '[[international journal of political economy'], ['hortscience'], ['europe-asia studies '], ['[[society for industrial and applied mathematics', 'siam review '], ['[[foreign policy analysis ', '[[oxford university press'], ['connections ', '[[partnership for peace consortium of defense academies and security studies institutes'], ['[[the university of chicago press', '[[the journal of modern history'], ['[[scientific american', 'scientific american'], ['[[canadian slavonic papers'], ['[[asian survey', '[[university of california press'], ['bmc public health '], ['[[the american historical review', '[[oxford university press'], ['journal for the study of religion'], ['[[slavic review', '[[cambridge university press'], ['family planning perspectives ', '[[guttmacher institute'], ['the review of politics '], ['the american slavic and east european review ', '[[association for slavic'], ['shs web of conferences '], ['[[foreign affairs'], ['the british medical journal '], ['[[slavic review'], ['[[the international history review', '[[taylor '], ['[[journal of the history of ideas', '[[university of pennsylvania press'], ['[[the american historical review', '[[oxford university press'], ['[[taylor ', '[[europe-asia studies'], ['[[university of pennsylvania press', '[[journal of the history of ideas'], ['[[the american mathematical monthly', '[[taylor '], ['[[review of central and east european law', '[[brill publishers'], ['[[war in history'], ['[[american political science association', '[[the american political science review'], ['[[canadian slavonic papers'], ['[[oxford university press', '[[journal of the american academy of religion'], ['[[the american historical review', '[[oxford university press'], ['[[quaternary international'], ['[[the monist', '[[oxford university press'], ['[[the russian review', '[[wiley '], ['[[journal of human evolution'], ['[[the russian review', '[[wiley '], ['[[journal of contemporary history'], ['[[raven'], ['[[comparative politics', 'comparative politics'], ['the [[university of chicago press', 'polity '], ['mayo clinic proceedings '], ['[[nature '], ['[[translation and literature', '[[edinburgh university press'], ['nature '], ['[[journal of the society of architectural historians'], ['[[russian history ', '[[brill publishers'], ['[[journal of multilingual and multicultural development', '[[european university institute'], ['[[geographical review', '[[taylor '], ['[[sage publishers', 'journal of modern european history ']]",78,32,0,146,0,12,177,0.1270358306188925,0.05211726384364821,0.23778501628664495,0.2785016286644951,0.0,0.4576547231270358,171,"['www.cia.gov', 'history.nasa.gov', 'www.cia.gov', 'www.cia.gov', 'www.nasa.gov', 'history.nasa.gov', 'nssdc.gsfc.nasa.gov', 'nssdc.gsfc.nasa.gov', 'solarsystem.nasa.gov', 'www.cia.gov', 'pubs.usgs.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'apps.fas.usda.gov', 'www.cia.gov', 'www.cia.gov', 'earthobservatory.nasa.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'rosstat.gov', 'www.cia.gov', 'crsreports.congress.gov', 'www.cia.gov', 'www.cia.gov', 'ac.gov', 'tourism.gov', 'www.loc.gov', 'www.historytoday.com', 'www.bbc.com', 'bp.com', 'www.britannica.com', 'www.britannica.com', 'www.britannica.com', 'www.nationalgeographic.com', 'www.uefa.com', 'www.bbc.com', 'www.bbc.com', 'thediplomat.com', 'www.nationalgeographic.com', 'www.bloomberg.com', 'www.theatlantic.com', 'www.economist.com', 'foreignpolicy.com', 'www.euractiv.com', 'www.theage.com', 'www.france24.com', 'www.trtworld.com', 'www.rbth.com', 'www.themoscowtimes.com', 'books.google.com', 'www.bbc.com', 'www.britannica.com', 'harvardpress.typepad.com', 'www.cnbc.com', 'books.google.com', 'www.expatica.com', 'www.bloomberg.com', 'www.wsj.com', 'www.fifa.com', 'books.google.com', 'www.aljazeera.com', 'knoema.com', 'www.themoscowtimes.com', 'www.economist.com', 'www.rbth.com', 'www.euronews.com', 'www.latimes.com', 'newzoo.com', 'www.bbc.com', 'www.bbc.com', 'www.merriam-webster.com', 'www.lingref.com', 'www.forbes.com', 'www.nytimes.com', 'kids.nationalgeographic.com', 'www.uefa.com', 'www.bloomberg.com', 'www.economist.com', 'books.google.com', 'www.newyorker.com', 'slate.com', 'www.britannica.com', 'tass.com', 'www.calvertjournal.com', 'docviewer.yandex.com', 'www.fifa.com', 'www.nytimes.com', 'www.newyorker.com', 'www.nytimes.com', 'researchfdi.com', 'www.nationalgeographic.com', 'qz.com', 'www.economy.com', 'books.google.com', 'www.themoscowtimes.com', 'www.nytimes.com', 'www.nationalgeographic.com', 'www.economist.com', 'www.washingtonpost.com', 'www.nytimes.com', 'www.washingtonpost.com', 'www.dw.com', 'www.bbc.com', 'www.historytoday.com', 'www.scientificamerican.com', 'www.scimagojr.com', 'books.google.com', 'books.google.com', 'www.dw.com', 'grantland.com', 'www.britannica.com', 'www.nationalgeographic.com', 'books.google.com', 'www.dw.com', 'www.usatoday.com', 'docviewer.yandex.com', 'www.wired.com', 'www.nytimes.com', 'www.britannica.com', 'www.nybooks.com', 'www.csmonitor.com', 'www.bbc.com', 'www.nytimes.com', 'www.britannica.com', 'www.latimes.com', 'www.vox.com', 'olympics.com', 'www.britannica.com', 'www.aa.com', 'thewest.com', 'www.themoscowtimes.com', 'www.britannica.com', 'www.voanews.com', 'www.topuniversities.com', 'www.ganintegrity.com', 'www.formula1.com', 'books.google.com', 'filmlinc.com', 'www.uefa.com', 'www.rbth.com', 'www.euronews.com', 'www.rbth.com', 'www.rbth.com', 'www.vox.com', 'www.nytimes.com', 'www.nytimes.com', 'www.voanews.com', 'www.dw.com', 'www.ft.com', 'www.straitstimes.com', 'www.rbth.com', 'books.google.com', 'www.discovermagazine.com', 'books.google.com', 'www.cnn.com', 'olympics.com', 'www.atlasobscura.com', 'www.atlasobscura.com', 'www.cbsnews.com', 'thediplomat.com', 'www.nytimes.com', 'edition.cnn.com', 'www.rbth.com', 'www.visualcapitalist.com', 'www.sbs.com', 'www.businessinsider.com', 'www.inverse.com', 'www.nytimes.com', 'www.themoscowtimes.com', 'www.britannica.com', 'www.bbc.com', 'books.google.com', 'www.themoscowtimes.com', 'imf.org', 'www.rferl.org', 'www.ucsusa.org', 'www.rferl.org', 'sgp.fas.org', 'www.rferl.org', 'www.armscontrol.org', 'www.ifri.org', 'www.amnesty.org', 'uis.unesco.org', 'www.rferl.org', 'www.irena.org', 'www.npr.org', 'ourworldindata.org', 'www.thearcticinstitute.org', 'rsf.org', 'library.oapen.org', 'worldroadstatistics.org', 'mjltm.org', 'sipri.org', 'data.worldbank.org', 'www.pbs.org', 'www.rand.org', 'www.irena.org', 'data.worldbank.org', 'sreda.org', 'globaldiplomacyindex.lowyinstitute.org', 'www.e-unwto.org', 'www.rferl.org', 'data.worldbank.org', 'www.pbs.org', 'www.rferl.org', 'data.worldbank.org', 'www.rferl.org', 'spectrum.ieee.org', 'files.stlouisfed.org', 'carnegieendowment.org', 'whc.unesco.org', 'power.lowyinstitute.org', 'www.hrw.org', 'www.rferl.org', 'unesdoc.unesco.org', 'data.worldbank.org', 'unesdoc.unesco.org', 'www.csen.org', 'www3.weforum.org', 'world-nuclear.org', 'www.unrisd.org', 'www.worldcat.org', 'daily.jstor.org', 'www.hrw.org', 'www.rferl.org', 'whc.unesco.org', 'www.bfi.org', 'data.worldbank.org', 'data.worldbank.org', 'www.paralympic.org', 'www.wilsoncenter.org', 'paleogeo.org', 'data.worldbank.org', 'www.unesco.org', 'hdr.undp.org', 'www.rferl.org', 'www.lowyinstitute.org', 'freedomhouse.org', 'education.rec.org', 'www.npr.org', 'data.worldbank.org', 'data.worldbank.org', 'www.nationalgeographic.org', 'www.transparency.org', 'www.jstor.org', 'worldenergy.org', 'unstats.un.org', 'education.rec.org', 'www.icrc.org', 'www.fao.org', 'www.iza.org', ['[[russian history '], ['[[cambridge university press', '[[slavic review'], ['politeja ', 'księgarnia akademicka '], ['[[the slavonic and east european review', '[[cambridge university press'], ['proceedings of the academy of political science ', '[[the academy of political science'], ['[[notes ', '[[music library association'], ['[[oxford university press', 'the musical quarterly'], ['[[parameters '], ['[[taylor ', '[[the international history review'], ['[[biographical memoirs of fellows of the royal society'], ['[[the american historical review', '[[oxford university press'], ['[[oecd'], ['[[sage publishing', '[[security dialogue'], ['[[oxford university press', 'oxford art journal'], ['the [[university of chicago press', '[[the quarterly review of biology'], ['[[nationalities papers'], ['[[slavic review', '[[cambridge university press'], ['[[oxford university press', '[[publius '], ['[[the slavonic and east european review', '[[modern humanities research association'], ['nature communications '], ['[[european journal of human genetics'], ['[[oxford university press', '[[the musical quarterly'], ['science '], ['[[the russian review'], ['the [[university of chicago press', '[[osiris'], ['[[the russian review', '[[wiley '], ['[[canadian international council', '[[sage publishing'], ['[[iranian studies', '[[taylor '], ['the world bank research observer ', '[[oxford university press'], ['caa ', '[[the art bulletin'], ['[[europe-asia studies'], ['[[college english', '[[national council of teachers of english'], ['[[council on foreign relations', '[[foreign affairs'], ['[[population and development review', '[[population council'], ['[[the russian review'], ['genomics ', '[[elsevier'], ['[[council on foreign relations', '[[foreign affairs'], ['[[academic studies press'], ['[[centre for european policy studies'], ['[[sage publishing', '[[social studies of science'], ['folklore'], ['[[royal historical society', '[[cambridge university press'], ['[[the russian review'], ['[[royal society', '[[obituary notices of fellows of the royal society'], [' [[nature '], ['[[journal of genocide research'], ['studies in conservation ', '[[taylor '], ['[[the russian review'], ['[[taylor ', '[[the american mathematical monthly'], ['[[third world quarterly', '[[taylor '], ['[[the journal of interdisciplinary history', 'the [[mit press'], ['[[journal of contemporary history', '[[sage publishing'], ['[[nationalities papers', '[[cambridge university press'], ['the art world'], ['[[notes '], ['[[princeton university', '[[contemporary european history'], ['the annals of the [[american academy of political and social science', '[[sage publishing'], ['rocky mountain modern language association ', 'rocky mountain review of language and literature'], ['journal of epidemiology and community health '], ['[[journal of world history', '[[university of hawaiʻi press'], ['[[european parliamentary research service', '[[european parliament'], ['[[russian history ', '[[brill publishers'], ['[[oxford university press', '[[journal of design history'], ['[[law ', '[[wiley '], ['[[taylor ', '[[europe-asia studies'], ['scientific data '], ['[[europe-asia studies', '[[taylor '], ['[[the russian review', '[[wiley '], ['[[academy of sciences of the soviet union', 'journal of the atmospheric sciences'], ['nature '], ['dance studies association ', '[[congress on research in dance'], ['[[university of california press', '[[asian survey'], ['communist and post-communist studies ', '[[university of california press'], ['the american political science review ', '[[american political science association'], [' [[the slavic and east european journal'], ['[[canadian slavonic papers'], ['[[perspectives on politics', '[[american political science association'], ['[[cambridge university press'], ['[[notes ', '[[music library association'], ['connections ', '[[partnership for peace consortium of defense academies and security studies institutes'], ['[[journal of economic perspectives', '[[harvard university'], ['[[brookings papers on economic activity', '[[brookings institution'], ['[[international organization', 'the [[mit press'], ['canadian medical association journal '], ['journal of innate immunity '], ['comparative politics ', '[[city university of new york'], ['[[annals of the association of american geographers', '[[taylor '], ['the soviet and post-soviet review', 'brill'], ['unwto world tourism barometer english version ', '[[world tourism organization'], ['[[university of pennsylvania press', '[[journal of the history of ideas'], ['alcohol and alcoholism '], ['[[the lancet'], ['geojournal '], ['[[nature photonics'], ['[[university of california press', '[[journal of the society of architectural historians'], ['[[nature photonics'], ['international journal on minority and group rights ', '[[brill publishers'], ['[[wiley ', '[[the russian review'], ['[[journal of contemporary history', '[[sage publishing'], ['[[the musical times'], ['nature '], ['[[brookings papers on economic activity'], ['[[journal of strategic security', '[[university of south florida'], ['[[the international history review'], ['[[past ', '[[oxford university press'], ['[[oxford university press', '[[music '], ['[[oecd'], ['[[europe-asia studies'], ['the journal of decorative and propaganda arts ', '[[florida international university'], ['[[the russian review', '[[wiley '], ['journal of international relations and development'], ['[[the johns hopkins university press', ' [[new literary history'], ['[[the russian review', '[[wiley '], ['[[international journal of environmental research and public health'], ['communist and post-communist studies', '[[university of california press'], ['[[university of california press', '[[chymia'], ['[[journal of contemporary history', '[[sage publishing'], ['[[the american political science review', '[[american political science association'], ['annual review of linguistics '], ['[[wiley ', '[[the russian review'], ['[[taylor ', '[[international journal of political economy'], ['hortscience'], ['europe-asia studies '], ['[[society for industrial and applied mathematics', 'siam review '], ['[[foreign policy analysis ', '[[oxford university press'], ['connections ', '[[partnership for peace consortium of defense academies and security studies institutes'], ['[[the university of chicago press', '[[the journal of modern history'], ['[[scientific american', 'scientific american'], ['[[canadian slavonic papers'], ['[[asian survey', '[[university of california press'], ['bmc public health '], ['[[the american historical review', '[[oxford university press'], ['journal for the study of religion'], ['[[slavic review', '[[cambridge university press'], ['family planning perspectives ', '[[guttmacher institute'], ['the review of politics '], ['the american slavic and east european review ', '[[association for slavic'], ['shs web of conferences '], ['[[foreign affairs'], ['the british medical journal '], ['[[slavic review'], ['[[the international history review', '[[taylor '], ['[[journal of the history of ideas', '[[university of pennsylvania press'], ['[[the american historical review', '[[oxford university press'], ['[[taylor ', '[[europe-asia studies'], ['[[university of pennsylvania press', '[[journal of the history of ideas'], ['[[the american mathematical monthly', '[[taylor '], ['[[review of central and east european law', '[[brill publishers'], ['[[war in history'], ['[[american political science association', '[[the american political science review'], ['[[canadian slavonic papers'], ['[[oxford university press', '[[journal of the american academy of religion'], ['[[the american historical review', '[[oxford university press'], ['[[quaternary international'], ['[[the monist', '[[oxford university press'], ['[[the russian review', '[[wiley '], ['[[journal of human evolution'], ['[[the russian review', '[[wiley '], ['[[journal of contemporary history'], ['[[raven'], ['[[comparative politics', 'comparative politics'], ['the [[university of chicago press', 'polity '], ['mayo clinic proceedings '], ['[[nature '], ['[[translation and literature', '[[edinburgh university press'], ['nature '], ['[[journal of the society of architectural historians'], ['[[russian history ', '[[brill publishers'], ['[[journal of multilingual and multicultural development', '[[european university institute'], ['[[geographical review', '[[taylor '], ['[[sage publishers', 'journal of modern european history ']]",25391,Require extended confirmed access (no expiry set),307576,31 October 2001,212.192.249.xxx ,21518,30,2001-10-31,2001-10,2001
138,138,Georgians,https://en.wikipedia.org/wiki/Georgians,69,2,"['10.1038/ejhg.2008.249', '10.3167/ame.2009.040205', '19107149', None, '2947100', None]","[['european journal of human genetics '], ['anthropology of the middle east']]",1,0,0,7,0,0,59,0.014492753623188406,0.0,0.10144927536231885,0.028985507246376812,0.0,0.043478260869565216,2,"['rbedrosian.com', 'books.google.com', 'books.google.com', 'books.google.com', 'rbedrosian.com', 'books.google.com', 'www.milliyet.com', 'www.iranicaonline.org', ['european journal of human genetics '], ['anthropology of the middle east']]",448609,Allow all users (no expiry set),36210,30 November 2003,80.191.134.142 ,3322,8,2003-11-30,2003-11,2003
139,139,North Macedonia,https://en.wikipedia.org/wiki/North_Macedonia,250,5,"['10.1038/s41467-020-19493-3', '10.1093/biosci/bix014', '10.4467/20834624sl.16.006.5152', '10.1016/j.sbspro.2012.05.001', '33293507', '28608869', None, None, '7723057', '5451287', None, None]","[['nature communications'], ['bioscience'], ['studia linguistica universitatis iagellonicae cracoviensis '], ['procedia - social and behavioral sciences']]",34,20,0,85,0,3,103,0.136,0.08,0.34,0.02,0.0,0.236,4,"['www.stat.gov', 'www.cia.gov', 'cia.gov', 'www.gov', 'www.stat.gov', 'macedonia.usaid.gov', 'makstat.stat.gov', 'www.stat.gov', 'www.instat.gov', 'stat.gov', 'www.stat.gov', 'www.stat.gov', 'www.moe.gov', 'www.stat.gov', 'www.mfa.gov', 'www.stat.gov', 'www.morm.gov', 'cia.gov', 'mfa.gov', 'www.stat.gov', 'books.google.com', 'idc-cema.com', 'www.slvesnik.com', 'books.google.com', 'www.kroraina.com', 'books.google.com', 'www.sbs.com', 'www.irishtimes.com', 'www.dnevnik.com', 'www.balkaneu.com', 'books.google.com', 'balkanalysis.com', 'books.google.com', 'www.bbc.com', 'books.google.com', 'www.mia.com', 'balkaninsight.com', 'media-2.web.britannica.com', 'balkaninsight.com', 'novinite.com', 'britannica.com', 'www.ft.com', 'books.google.com', 'books.google.com', 'nuwireinvestor.com', 'foreignpolicy.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'www.dw.com', 'www.beinsports.com', 'nationalpost.com', 'kroraina.com', 'books.google.com', 'www.bbc.com', 'books.google.com', 'euractiv.com', 'www.reuters.com', 'books.google.com', 'balkaninsight.com', 'www.britannica.com', 'www.etymonline.com', 'books.google.com', 'www.ethnologue.com', 'books.google.com', 'slate.com', 'books.google.com', 'books.google.com', 'www.dw.com', 'www.findarticles.com', 'www.balkaninsight.com', 'www.setimes.com', 'balkaninsight.com', 'euratlas.com', 'thestar.com', 'books.google.com', 'britannica.com', 'www.bbc.com', 'www.balkaninsight.com', 'books.google.com', 'books.google.com', 'www.cp24.com', 'www.kroraina.com', 'www.euractiv.com', 'books.google.com', 'www.dw.com', 'books.google.com', 'www.euronews.com', 'books.google.com', 'www.novinite.com', 'www.britannica.com', 'britannica.com', 'www.aljazeera.com', 'www.dw.com', 'books.google.com', 'books.google.com', 'makstack.com', 'www.reuters.com', 'www.reuters.com', 'novinite.com', 'www.dw.com', 'uefa.com', 'www.reuters.com', 'www.findarticles.com', 'books.google.com', 'promacedonia.org', 'www.ushmm.org', 'www.un.org', 'www.pewforum.org', 'rsf.org', 'heritage.org', 'dergipark.org', 'doingbusiness.org', 'devdata.worldbank.org', 'www.un.org', 'www.rferl.org', 'lnweb90.worldbank.org', 'www.oic.org', 'europeandcis.undp.org', 'www.ejil.org', 'visionofhumanity.org', 'worldbank.org', 'www.rferl.org', 'www.promacedonia.org', 'www.rferl.org', 'greekembassy.org', 'www.livius.org', 'sr.wikisource.org', 'hdr.undp.org', 'sr.wikisource.org', 'www.imf.org', 'transparency.org', 'www.un.org', 'www.ushmm.org', 'www.hrw.org', 'hdr.undp.org', 'www.worldbank.org', 'www.un.org', 'web.amnesty.org', ['nature communications'], ['bioscience'], ['studia linguistica universitatis iagellonicae cracoviensis '], ['procedia - social and behavioral sciences']]",23564616,Require administrator access (no expiry set),178677,26 February 2002,195.170.0.24 ,10404,15,2002-02-26,2002-02,2002
140,140,Montenegro,https://en.wikipedia.org/wiki/Montenegro,135,2,"['10.1093/biosci/bix014', '10.1038/s41467-020-19493-3', '28608869', '33293507', '5451287', '7723057']","[['bioscience'], ['nature communications']]",29,7,0,53,0,1,44,0.21481481481481482,0.05185185185185185,0.3925925925925926,0.014814814814814815,0.0,0.2814814814814815,2,"['www.ttk.gov', 'www.gov', 'mvpei.gov', 'www.gov', 'www.cia.gov', 'mvp.gov', '2009-2017.state.gov', 'books.google.com', 'www.myguidemontenegro.com', 'balkaninsight.com', 'www.reuters.com', 'books.google.com', 'in.reuters.com', 'www.bbc.com', 'www.irishtimes.com', 'www.lonelyplanet.com', 'adventureworldmagazineonline.com', 'abcnews.go.com', 'books.google.com', 'abcnews.go.com', 'www.myguidemontenegro.com', 'www.euronews.com', 'www.nytimes.com', 'www.bbc.com', 'books.google.com', 'www.washingtontimes.com', 'visit-montenegro.com', 'blogs.nationalgeographic.com', 'www.balkaninsight.com', 'www.ft.com', 'www.todayszaman.com', 'www.britannica.com', 'www.jamesbondlifestyle.com', 'total-waterpolo.com', 'books.google.com', 'kotoronline.com', 'europeanwesternbalkans.com', 'www.montenegro.com', 'europeanwesternbalkans.com', 'sfmission.com', 'www.bbc.com', 'www.wsj.com', 'www.dw.com', 'books.google.com', 'croatiatraveller.com', 'sonypictures.com', 'books.google.com', 'www.balkans.com', 'www.nytimes.com', 'www.foreignpolicyjournal.com', 'books.google.com', 'www.nytimes.com', 'rs.n1info.com', 'www.visit-montenegro.com', 'www.wsj.com', 'travel.yahoo.com', 'books.google.com', 'www.aljazeera.com', 'rs.n1info.com', 'www.voanews.com', 'monstat.org', 'yihr.org', 'hosted.ap.org', 'www.rferl.org', 'www.un.org', 'www.nationsonline.org', 'freedomhouse.org', 'hdr.undp.org', 'gutenberg.org', 'montenegro.org', 'hosted.ap.org', 'www.jstor.org', 'imf.org', 'www.rferl.org', 'freedomhouse.org', 'www.occrp.org', 'www.iso.org', 'www.monstat.org', 'www.heritage.org', 'aceproject.org', 'hdr.undp.org', 'imf.org', 'www.monstat.org', 'www.monstat.org', 'www.slobodnaevropa.org', 'www.monstat.org', 'njegos.org', 'www.slobodnaevropa.org', 'devdata.worldbank.org', ['bioscience'], ['nature communications']]",20760,Require administrator access (no expiry set),119801,16 December 2001,David Parker ,9674,41,2001-12-16,2001-12,2001
141,141,Czech Republic,https://en.wikipedia.org/wiki/Czech_Republic,232,10,"['10.1111/j.1467-9515.2009.00654.x', '10.1002/ijop.12607', '10.1093/past/153.1.164', '10.1093/biosci/bix014', '10.1038/s41467-020-19493-3', '10.1175/mwr-d-15-0298.1', '10.1007/s00704-018-2553-y', '10.1093/oep/gpt036', '10.5334/ijic.8', '10.1515/bjlp-2015-0004', None, '31304980', None, '28608869', '33293507', None, None, None, '16902697', None, None, None, None, '5451287', '7723057', None, None, None, '1534002', None]","[['social policy '], ['international journal of psychology '], ['past and present'], ['bioscience'], ['nature communications'], [' mon. wea. rev. '], [' theor. appl. climatol. '], ['oxford economic papers'], ['int j integr care '], ['baltic journal of law ']]",28,7,0,60,0,1,127,0.1206896551724138,0.03017241379310345,0.25862068965517243,0.04310344827586207,0.0,0.1939655172413793,10,"['travel.state.gov', '2009-2017.state.gov', 'www.cia.gov', 'cia.gov', 'www.cia.gov', 'www.portal.gov', 'www.cia.gov', 'www.czech-research.com', 'articles.latimes.com', 'www.nytimes.com', 'groups.yahoo.com', 'books.google.com', 'www.economist.com', 'books.google.com', 'thenextweb.com', 'www.collinsdictionary.com', 'blog.euromonitor.com', 'books.google.com', 'wingia.com', 'travelguidepro.com', 'books.google.com', 'www.czechia-initiative.com', 'www.amazon.com', 'www.henleyglobal.com', 'news.com', 'www.wingia.com', 'www.bleepingcomputer.com', 'www.kftv.com', 'books.google.com', 'www.oed.com', 'books.google.com', 'factsmaps.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'www.sciencefriday.com', 'www.huffingtonpost.com', 'www.reuters.com', 'books.google.com', 'books.google.com', 'www.scimagoir.com', 'www.allianz.com', 'books.google.com', 'www.skoda-storyboard.com', 'www.britannica.com', 'healthpowerhouse.com', 'www.dw.com', 'www.ft.com', 'www.myczechrepublic.com', 'www.bbc.com', 'ahdictionary.com', 'books.google.com', 'www.usnews.com', 'www.yeyeagency.com', 'www.czechtourism.com', 'dw.com', 'www.openculture.com', 'www.praguepost.com', 'books.google.com', 'en.oxforddictionaries.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.praguepost.com', 'www.czechinvest.org', 'imf.org', 'nobelprize.org', 'unesco.org', 'hdr.undp.org', 'web.worldbank.org', 'ushmm.org', 'unstats.un.org', 'www.jewishvirtuallibrary.org', 'www.pewforum.org', 'imf.org', 'reports.weforum.org', 'oecd.org', 'svu2000.org', 'www.worldcat.org', 'www.museeprotestant.org', 'www.heritage.org', 'www.globalinnovationindex.org', 'visionofhumanity.org', 'imf.org', 'undp.org', 'whc.unesco.org', 'unterm.un.org', 'www.wilsoncenter.org', 'www.worldjewishcongress.org', 'rsf.org', 'hdr.undp.org', 'reports.weforum.org', ['social policy '], ['international journal of psychology '], ['past and present'], ['bioscience'], ['nature communications'], [' mon. wea. rev. '], [' theor. appl. climatol. '], ['oxford economic papers'], ['int j integr care '], ['baltic journal of law ']]",5321,Require administrator access (no expiry set),169281,20 July 2001,Koyaanis Qatsi ,10524,13,2001-07-20,2001-07,2001
142,142,Culture of Telangana,https://en.wikipedia.org/wiki/Culture_of_Telangana,50,1,"['10.1080/02666030.1993.9628458', None, None]",[['south asian studies']],3,6,0,31,0,0,9,0.06,0.12,0.62,0.02,0.0,0.2,1,"['www.telangana.gov', 'ccrtindia.gov', 'aptdc.gov', 'cbfcindia.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'timesofindia.indiatimes.com', 'indianexpress.com', 'www.thehindu.com', 'www.britannica.com', 'deccanchronicle.com', 'www.hindu.com', 'www.thehindu.com', 'www.siasat.com', 'articles.timesofindia.indiatimes.com', 'travel.outlookindia.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'www.info4india.com', 'www.indiainfoweb.com', 'www.thehindu.com', 'www.languageinindia.com', 'www.hindu.com', 'books.google.com', 'www.hindu.com', 'www.hindu.com', 'www.indiayogi.com', 'guinnessworldrecords.com', 'books.google.com', 'travel.cnn.com', 'www.astroved.com', 'www.thehindu.com', 'www.hindu.com', 'www.thehindu.com', 'gizmodo.com', 'timesofindia.indiatimes.com', 'stjohnschurchcsi.org', 'vemulawadatemple.org', 'bhadrachalarama.org', ['south asian studies']]",43345266,Allow all users (no expiry set),41804,19 July 2014,Hariehkr ,334,0,2014-07-19,2014-07,2014
143,143,Kongu Nadu,https://en.wikipedia.org/wiki/Kongu_Nadu,63,0,[],[],2,0,0,41,0,0,20,0.031746031746031744,0.0,0.6507936507936508,0.0,0.0,0.031746031746031744,0,"['papers.ssrn.com', 'www.krepublishers.com', 'www.business-standard.com', 'www.thehindu.com', 'www.thehindu.com', 'www.hindu.com', 'www.hindu.com', 'www.hindu.com', 'www.rediff.com', 'www.hinduonnet.com', 'www.news18.com', 'www.hindu.com', 'www.hindu.com', 'books.google.com', 'www.hindu.com', 'articles.timesofindia.indiatimes.com', 'www.thehindubusinessline.com', 'tamilartsacademy.com', 'books.google.com', 'www.bbc.com', 'timesofindia.indiatimes.com', 'www.thenewsminute.com', 'www.britannica.com', 'www.thehindu.com', 'www.newindianexpress.com', 'www.iskconhighertaste.com', 'www.thequint.com', 'books.google.com', 'hindu.com', 'www.hindu.com', 'www.hindu.com', 'www.newindianexpress.com', 'www.thehindu.com', 'books.google.com', 'www.hindustantimes.com', 'www.news18.com', 'www.thehindu.com', 'tamil.abplive.com', 'www.livemint.com', 'www.thehindu.com', 'www.indiatimes.com', 'www.jstor.org', 'apmn.icimod.org']",1937921,Allow all users (no expiry set),36896,25 May 2005,Tom Radulovich ,2392,7,2005-05-25,2005-05,2005
144,144,Pastirma,https://en.wikipedia.org/wiki/Pastirma,52,9,"['10.2307/632150', '10.1016/j.jef.2018.02.004', '10.1093/acref/9780192806819.001.0001', '10.1016/j.lwt.2009.05.016', '10.1016/j.meatsci.2006.04.001', '10.1525/ctx.2007.6.3.67', '10.1016/j.foodres.2017.09.094', '10.1016/b978-0-12-384731-7.00197-5', '10.1016/j.meatsci.2013.03.021', None, None, None, None, '22062846', None, '29195938', None, '23608196', None, None, None, None, None, None, None, None, None]","[[' the journal of hellenic studies'], [' journal of ethnic foods'], [' oxford university press'], [' lwt - food science and technology'], [' meat science'], [' contexts'], [' food research international'], ['elsevier'], [' meat science']]",0,0,0,31,0,0,12,0.0,0.0,0.5961538461538461,0.17307692307692307,0.0,0.17307692307692307,9,"['www.youtube.com', 'books.google.com', 'www.youtube.com', 'armenianweekly.com', 'books.google.com', 'books.google.com', 'www.youtube.com', 'www.youtube.com', 'www.youtube.com', 'books.google.com', 'books.google.com', 'www.youtube.com', 'www.youtube.com', 'books.google.com', 'www.youtube.com', 'www.youtube.com', 'www.youtube.com', 'books.google.com', 'www.youtube.com', 'books.google.com', 'books.google.com', 'www.youtube.com', 'books.google.com', 'www.youtube.com', 'thisweekinpalestine.com', 'www.youtube.com', 'www.cumhuriyet.com', 'www.sabah.com', 'books.google.com', 'articles.latimes.com', 'books.google.com', [' the journal of hellenic studies'], [' journal of ethnic foods'], [' oxford university press'], [' lwt - food science and technology'], [' meat science'], [' contexts'], [' food research international'], ['elsevier'], [' meat science']]",1226536,Allow all users (no expiry set),25370,30 November 2004,85.96.11.162 ,893,0,2004-11-30,2004-11,2004
145,145,Laz people,https://en.wikipedia.org/wiki/Laz_people,67,3,"['10.1080/00263206.2011.652778', '10.1163/ej.9789004163089.i-1122.306', '10.7256/1994-1471.2014.5.9758', None, None, None, None, None, None]","[['middle eastern studies'], ['brill'], ['актуальные проблемы российского права']]",8,2,0,15,0,0,39,0.11940298507462686,0.029850746268656716,0.22388059701492538,0.04477611940298507,0.0,0.19402985074626866,3,"['dspace.nplg.gov', 'nplg.gov', 'books.google.com', 'www.hurriyetdailynews.com', 'www.languagesandnumbers.com', 'www.ethnologue.com', 'www.britannica.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.yeniansiklopedi.com', 'www.ethnologue.com', 'referenceworks.brillonline.com', 'www.ethnologue.com', 'www.dailysabah.com', 'encyclopedia.com', 'i-cias.com', 'lazca.org', 'www.bianet.org', 'chai-khana.org', 'newadvent.org', 'www.usefoundation.org', 'www.unesco.org', 'www.wdl.org', 'usefoundation.org', ['middle eastern studies'], ['brill'], ['актуальные проблемы российского права']]",5497767,Require autoconfirmed or confirmed access (no expiry set),50904,9 June 2006,Khoikhoi ,948,0,2006-06-09,2006-06,2006
146,146,Iran,https://en.wikipedia.org/wiki/Iran,572,7,"['10.1017/s0017816000007926', '10.1007/bf00161055', '10.1353/pew.2002.0030', '10.1002/jtr.862', '10.1017/s0035869x0012965x', '10.1080/10163270802006321', '10.1038/s41467-020-19493-3', None, None, None, None, None, None, '33293507', None, None, None, None, None, None, '7723057']","[['the harvard theological review'], ['indo-iranian journal ', 'brill '], ['philosophy east and west ', 'university of hawai'], ['international journal of tourism research'], [' journal of the royal asiatic society of great britain '], [' korean journal of defense analysis'], ['nature communications']]",91,14,0,305,0,10,146,0.1590909090909091,0.024475524475524476,0.5332167832167832,0.012237762237762238,0.0,0.1958041958041958,7,"['cia.gov', 'www.cia.gov', 'cia.gov', 'eia.doe.gov', 'www.state.gov', 'www.loc.gov', 'www.uktradeinvest.gov', 'www.cia.gov', 'www.mfa.gov', 'lcweb2.loc.gov', 'www.state.gov', 'www.justice.gov', 'www.usgs.gov', 'webarchive.loc.gov', 'www.bbc.com', 'iran-daily.com', 'books.google.com', 'ivarta.com', 'www.timesofisrael.com', 'books.google.com', 'www.al-monitor.com', 'books.google.com', 'www.iranchamber.com', 'www.findarticles.com', 'www.studentpulse.com', 'www.reuters.com', 'pronounce.voanews.com', 'al-monitor.com', 'www2.irna.com', 'pbase.com', 'sports.espn.go.com', 'arabiancampus.com', 'www.eiu.com', 'massoudmehrabi.com', 'www.tabletmag.com', 'books.google.com', 'www.religionfacts.com', 'books.google.com', 'apnews.com', 'books.google.com', 'articles.latimes.com', 'abc-of-mountaineering.com', 'books.google.com', 'www.washingtonpost.com', 'chicagotribune.com', 'www.nytimes.com', 'books.google.com', 'www.thenewsminute.com', 'books.google.com', 'www.mysteryofiran.com', 'payvand.com', 'www.ancientscripts.com', 'www.al-monitor.com', 'thediplomat.com', 'books.google.com', 'theheritagetrust.wordpress.com', 'www.nytimes.com', 'www.britannica.com', 'www.tehrantimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'historic-uk.com', 'books.google.com', 'books.google.com', 'payvand.com', 'www.nanovip.com', 'financialtribune.com', 'www.scimagolab.com', 'books.google.com', 'destinationiran.com', 'books.google.com', 'books.google.com', 'www.reuters.com', 'www.nbcnews.com', 'www.nybooks.com', 'books.google.com', 'books.google.com', 'www.reuters.com', 'books.google.com', 'kayhanlife.com', 'www.reuters.com', 'books.google.com', 'www.al-monitor.com', 'www.britannica.com', 'news.xinhuanet.com', 'www.aljazeera.com', 'books.google.com', 'www.nytimes.com', 'www.washingtonpost.com', 'books.google.com', 'www.france24.com', 'books.google.com', 'www.nytimes.com', 'boioks.google.com', 'www.thedailybeast.com', 'parstimes.com', 'www.newsweek.com', 'books.google.com', 'www.tehrantimes.com', 'books.google.com', 'encarta.msn.com', 'www.bbc.com', 'destinationiran.com', 'observers.france24.com', 'books.google.com', 'news.yahoo.com', 'www.haaretz.com', 'www.nytimes.com', 'books.google.com', 'books.google.com', 'iranwire.com', 'www.payvand.com', 'www.persiansarenotarabs.com', 'observers.france24.com', 'www.iran-daily.com', 'billypenn.com', 'polomuseum.com', 'books.google.com', 'financialtribune.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'azargoshnasp.com', 'ahdictionary.tumblr.com', 'www.reuters.com', 'america.aljazeera.com', 'www.wsj.com', 'en.mehrnews.com', 'www.payvand.com', 'sacredsites.com', 'www.cnn.com', 'animation-festivals.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.tasnimnews.com', 'books.google.com', 'iranchamber.com', 'books.google.com', 'iranintl.com', 'www.reuters.com', 'www.britannica.com', 'www.tehrantimes.com', 'www.britannica.com', 'www.radiofarda.com', 'www.iran-daily.com', 'books.google.com', 'books.google.com', 'www.turquoisepartners.com', 'www.thebusinessyear.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'iranchamber.com', 'www.merriam-webster.com', 'www.bernama.com', 'old.iran-daily.com', 'archaeology.about.com', 'books.google.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.al-monitor.com', 'www.iran-daily.com', 'payvand.com', 'books.google.com', 'www.dw.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.britannica.com', 'www.internetworldstats.com', 'books.google.com', 'payvand.com', 'books.google.com', 'washingtonjewishweek.com', 'www.alexa.com', 'iranchamber.com', 'aa.com', 'books.google.com', 'www.iranian.com', 'www.bbc.com', 'www.economist.com', 'www.timesofisrael.com', 'books.google.com', 'books.google.com', 'usatoday30.usatoday.com', 'payvand.com', 'www.britannica.com', 'www.britannica.com', 'books.google.com', 'www.foxnews.com', 'heraldextra.com', 'books.google.com', 'books.google.com', 'news.yahoo.com', 'transoxiana.com', 'www.nbcnews.com', 'worldpopulationreview.com', 'www.nytimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'britannica.com', 'books.google.com', 'www.thebaghdadpost.com', 'bbcpersian.com', 'books.google.com', 'books.google.com', 'smithsonianmag.com', 'books.google.com', 'books.google.com', 'allaboutturkey.com', 'books.google.com', 'www.theatlantic.com', 'books.google.com', 'levity.com', 'dw.com', 'www.iran-daily.com', 'www.iran-daily.com', 'books.google.com', 'books.google.com', 'fifa.com', 'books.google.com', 'photius.com', 'fsmitha.com', 'aipsmedia.com', 'www.sfgate.com', 'books.google.com', 'books.google.com', 'www.ft.com', 'www.newsweek.com', 'books.google.com', 'iran-daily.com', 'news.xinhuanet.com', 'books.google.com', 'traveldocs.com', 'books.google.com', 'www.stalbertgazette.com', 'payvand.com', 'books.google.com', 'www.payvand.com', 'www.economist.com', 'www.realmofhistory.com', 'payvand.com', 'books.google.com', 'middle-east-online.com', 'www.iranchamber.com', 'www.hollandsentinel.com', 'www.washingtonpost.com', 'en.allexperts.com', 'foreignpolicy.com', 'www.britannica.com', 'rockclimbing.com', 'www.aljazeera.com', 'books.google.com', 'computerworld.com', 'encarta.msn.com', 'washingtontimes.com', 'english.aawsat.com', 'snowseasoncentral.com', 'books.google.com', 'oilprice.com', 'books.google.com', 'www.reuters.com', 'books.google.com', 'www.slate.com', 'books.google.com', 'english.aawsat.com', 'books.google.com', 'worldofvolley.com', 'panshin.com', 'iranchamber.com', 'books.google.com', 'www.iran-daily.com', 'books.google.com', 'books.google.com', 'theconversation.com', 'books.google.com', 'art-arena.com', 'farsnews.com', 'books.google.com', 'www.google.com', 'en.numista.com', 'financialtribune.com', 'books.google.com', 'books.google.com', 'books.google.com', 'occawlonline.pearsoned.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'money.cnn.com', 'books.google.com', 'books.google.com', 'iran-daily.com', 'iranonline.com', 'www.trtworld.com', 'wsj.com', 'boioks.google.com', 'www.stalbertgazette.com', 'www.al-monitor.com', 'www.nbcnews.com', '(www.dw.com', 'books.google.com', 'observers.france24.com', 'www.guinnessworldrecords.com', 'books.google.com', 'weather-and-climate.com', 'en.oxforddictionaries.com', 'www.iran-daily.com', 'observers.france24.com', 'books.google.com', 'info.worldbank.org', 'www.hrw.org', 'www.c-span.org', 'www.iranicaonline.org', 'www.iranicaonline.org', 'www.iucnredlist.org', 'www.iranicaonline.org', 'esa.un.org', 'www.hamsaweb.org', 'uis.unesco.org', 'www.amar.org', 'faostat.fao.org', 'wes.org', 'www.iranicaonline.org', 'www.un.org', 'irinnews.org', 'www.iranicaonline.org', 'www.criticalthreats.org', 'www.hrw.org', 'www.amnesty.org', 'stats.oecd.org', 'washingtoninstitute.org', 'www.worldaffairsjournal.org', 'www.hrw.org', 'www.globalsecurity.org', 'data.worldbank.org', 'www.iranicaonline.org', 'imf.org', 'pbs.org', 'data.worldbank.org', 'www.un.org', 'www.iranicaonline.org', 'www.iranicaonline.org', 'data.worldbank.org', 'migrationinformation.org', 'rsf.org', 'www.iranicaonline.org', 'www.iranicaonline.org', 'ancawr.org', 'faostat3.fao.org', 'stats.uis.unesco.org', 'www.amnesty.org', 'www.amnesty.org', 'www.iranicaonline.org', 'www.iranhrdc.org', 'www.iranicaonline.org', 'www.amar.org', 'www.iranicaonline.org', 'whc.unesco.org', 'www.worldvaluessurvey.org', 'www.iranicaonline.org', 'freedomhouse.org', 'iranicaonline.org', 'ourworldindata.org', 'www.unesco.org', 'iranicaonline.org', 'data.worldbank.org', 'www.globalsecurity.org', 'unesco.org', 'fa.wikisource.org', 'www.jstor.org', 'www.iranicaonline.org', 'www.iranicaonline.org', 'isg-mit.org', 'treaties.un.org', 'globalsecurity.org', 'iran-shutdown.amnesty.org', 'www.amar.org', 'www.iranicaonline.org', 'ourworldindata.org', 'www.britishmuseum.org', 'www.rferl.org', 'gamaan.org', 'www.iranicaonline.org', 'www.gloria-center.org', 'unesco.org', 'www.rferl.org', 'electionguide.org', 'www.unhcr.org', 'www.iranicaonline.org', 'www.sci.org', 'globalsecurity.org', 'rsf.org', 'hdr.undp.org', 'go.worldbank.org', 'www.washingtoninstitute.org', 'undocs.org', 'www.eurasianhome.org', 'www.fidh.org', 'www.iranicaonline.org', 'www.iranicaonline.org', ['the harvard theological review'], ['indo-iranian journal ', 'brill '], ['philosophy east and west ', 'university of hawai'], ['international journal of tourism research'], [' journal of the royal asiatic society of great britain '], [' korean journal of defense analysis'], ['nature communications']]",14653,Require administrator access (no expiry set),318320,22 October 2001,Zundark ,20086,25,2001-10-22,2001-10,2001
147,147,Mexico,https://en.wikipedia.org/wiki/Mexico,478,15,"['10.1215/00182168-36.3.309', '10.1353/jaas.2011.0029', '10.1017/s0022216x00017533', '10.1017/s026021051000135x', '10.18111/9789284419029', '10.1353/tam.2001.0109', '10.1525/mex.2015.31.2.218', '10.1146/annurev.anthro.26.1.129', '10.1007/s12394-010-0074-7', '10.1590/s0036-36342011000200005', '10.1177/0003122410378232', '10.29043/liminar.v6i1.263', '10.1016/s0277-9536(97)00023-3', '10.1038/s41467-020-19493-3', None, None, None, None, None, None, None, None, None, '21537803', None, None, '9381229', '33293507', None, None, None, None, None, None, None, None, None, None, None, None, None, '7723057']","[['hispanic american historical review '], ['journal of asian american studies'], [' journal of latin american studies '], ['review of international studies '], ['world tourism organization '], ['the americas', 'university of utah press'], ['mexican studies'], ['annual review of anthropology '], [' identity in the information society'], ['salud pública de méxico '], ['american sociological review ', 'american sociological association '], ['liminar '], ['social science '], ['nature communications ']]",89,18,0,173,0,2,181,0.18619246861924685,0.03765690376569038,0.3619246861924686,0.03138075313807531,0.0,0.25523012552301255,14,"['www.cia.gov', 'www.cia.gov', 'factfinder.census.gov', 'www.cia.gov', '2001-2009.state.gov', 'www.cia.gov', 'www.cia.gov', 'www.eia.doe.gov', 'www.cia.gov', 'cia.gov', 'www.cia.gov', 'state.gov', 'travel.state.gov', 'www.cia.gov', 'eia.doe.gov', 'www.ustreas.gov', 'www.dea.gov', 'www.loc.gov', 'books.google.com', 'azcentral.com', 'www.latinobookreview.com', 'www.milenio.com', 'books.google.com', 'photius.com', 'www.britannica.com', 'themazatlanpost.com', 'eleconomista.com', 'www.sandiegometro.com', 'www.bbvaresearch.com', 'books.google.com', 'guadalajarareporter.com', 'books.google.com', 'www.ft.com', 'www.sipuebla.com', 'mapscaping.com', 'www.milenio.com', 'www.emayzine.com', 'www.eluniversal.com', 'www.sfgate.com', 'www.mediotiempo.com', 'books.google.com', 'online.wsj.com', 'www.esmas.com', 'www.bloomberg.com', 'www.aicm.com', 'www.huffpost.com', 'www.milenio.com', 'www.latimes.com', 'charroazteca.com', 'www.rsssf.com', 'www.clutejournals.com', 'books.google.com', 'books.google.com', 'mexiconewsdaily.com', 'www.americaeconomia.com', 'pacificallianceblog.com', 'impreso.milenio.com', 'www.eleconomista.com', 'edition.cnn.com', 'www.ft.com', 'mexico.as.com', 'www.vallartadaily.com', 'www.britannica.com', 'www.elsoldemexico.com', 'www.jornada.com', 'books.google.com', 'www.dina.com', 'www.forbes.com', 'www.bbc.com', 'www.todaytranslations.com', 'somosprimos.com', 'spaceref.com', 'latinola.com', 'expatforum.com', 'www.photius.com', 'articlealley.com', 'books.google.com', 'www.marca.com', 'www.elfinanciero.com', 'www.jornada.com', 'www.economist.com', 'www.forbes.com', 'www.tlahui.com', 'books.google.com', 'books.google.com', 'www.concacaf.com', 'cnnsi.com', 'money.cnn.com', 'books.google.com', 'books.google.com', 'www.washingtonpost.com', 'prnewswire.com', 'globerove.com', 'www.nytimes.com', 'icabo.com', 'www.oxanstore.com', 'www.accessmylibrary.com', 'upi.com', 'tech.com', 'www.rigzone.com', 'www.elfinanciero.com', 'www.mediotiempo.com', 'www.nbcnews.com', 'books.google.com', 'www.autoblog.com', 'www.britannica.com', 'cervantesvirtual.com', 'insearchoflostplaces.com', 'www.satmex.com', 'www.liquor.com', 'terra.com', 'www.britannica.com', 'loutardeliberee.com', 'www.aicm.com', 'www.eluniversal.com', 'books.google.com', 'noticieros.televisa.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.mb.com', 'books.google.com', 'books.google.com', 'www.washingtonpost.com', 'www.fiba.com', 'www.britannica.com', 'www.nytimes.com', 'www.britannica.com', 'www.bbc.com', 'www.forbes.com', 'www.inside-mexico.com', 'www.grammarly.com', 'www.catholicnewsagency.com', 'books.google.com', 'thediplomat.com', 'www.systra.com', 'azcentral.com', 'www.budde.com', 'theconversation.com', 'elpais.com', 'books.google.com', 'books.google.com', 'www.oxanstore.com', 'www.investopedia.com', 'www.latinobookreview.com', 'www.rsssf.com', 'books.google.com', 'britannica.com', 'www.chemicool.com', 'www.iie.com', 'www.eluniversal.com', 'www.washingtontimes.com', 'www.cityexpress.com', 'books.google.com', 'www.thoughtco.com', 'books.google.com', 'www.economist.com', 'www.nytimes.com', 'www.huffingtonpost.com', 'www.reuters.com', 'books.google.com', 'www.autoexplora.com', 'www.pwc.com', 'snellwilcox.com', 'www.scmp.com', 'books.google.com', 'adherents.com', 'articles.latimes.com', 'books.google.com', 'www.iie.com', 'www.nytimes.com', 'mapscaping.com', 'busquedas.gruporeforma.com', 'www.arqhys.com', 'www.americaeconomia.com', 'foreignpolicy.com', 'www.milenio.com', 'www.elsoldemexico.com', 'www.britannica.com', 'www.mexicoescultura.com', 'www.dineroenimagen.com', 'books.google.com', 'books.google.com', 'www.lapatilla.com', 'www.milenio.com', 'lasillarota.com', 'www.stratfor.com', 'www.cronica.com', 'www.eluniversal.com', 'ancientcivilizationsworld.com', 'www.oecd-ilibrary.org', 'www.newadvent.org', 'oregon.conevyt.org', 'www.worldcat.org', 'www.globalsecurity.org', 'www.insightcrime.org', 'www.oecd.org', 'www.inegi.org', 'www.scielo.org', 'www.oecd.org', 'dallasfed.org', 'www.oecd.org', 'michaeljournal.org', 'www.pri.org', 'www.inegi.org', 'www.inegi.org', 'www.foreignaffairs.org', 'ierd.prd.org', 'www.conapred.org', 'www.conapred.org', 'nobelprize.org', 'report.globalintegrity.org', 'www.cfr.org', 'stats.oecd.org', 'www.prd.org', 'hdr.undp.org', 'www.koreauspartnership.org', 'www.theworldwar.org', 'www.beta.inegi.org', 'www.pen.org', 'www.cambridge.org', 'www.donquijote.org', 'ei.britishcouncil.org', 'diplomaticosescritores.org', 'www.odca.org', 'mx.ambafrance.org', 'www.fundacionunam.org', 'www.un.org', 'www.overseasvotefoundation.org', 'www.inegi.org', 'www.migrationpolicy.org', 'www.francophonie.org', 'www.npr.org', 'visionofhumanity.org', 'wayback.archive-it.org', 'opanal.org', 'hdr.undp.org', 'normateca.ife.org', 'www.inegi.org', 'www3.inegi.org', 'whc.unesco.org', 'www.aguas.org', 'theglobalamericans.org', 'www.inegi.org', 'www.un.org', 'siteresources.worldbank.org', 'www.cambridge.org', 'redalyc.org', 'www.femexfut.org', 'normateca.ife.org', 'www.conapred.org', 'newsroom.lds.org', 'www.inegi.org', 'www.scielo.org', 'www.latinamericanstudies.org', 'siteresources.worldbank.org', 'mexicka.org', 'data.oecd.org', 'agua.org', 'oxfamblogs.org', 'normateca.ife.org', 'whc.unesco.org', 'thecatalist.org', 'www.imf.org', 'opanal.org', 'aleph.org', 'wayback.archive-it.org', 'www.imef.org', 'www.eclac.org', 'www.catholic.org', 'www.pbs.org', 'www.globalpolicy.org', 'cuentame.inegi.org', 'www.sciencemag.org', 'www2.ohchr.org', 'www3.weforum.org', 'treaties.un.org', 'fas.org', 'lopezobrador.org', ['hispanic american historical review '], ['journal of asian american studies'], [' journal of latin american studies '], ['review of international studies '], ['world tourism organization '], ['the americas', 'university of utah press'], ['mexican studies'], ['annual review of anthropology '], [' identity in the information society'], ['salud pública de méxico '], ['american sociological review ', 'american sociological association '], ['liminar '], ['social science '], ['nature communications ']]",3966054,Require extended confirmed access (no expiry set),319104,13 August 2002,Brion VIBBER ,15851,144,2002-08-13,2002-08,2002
148,148,Wales,https://en.wikipedia.org/wiki/Wales,430,1,"['10.1144/gsl.jgs.1852.008.01-02.20', None, None]",[['q. j. geol. soc. lond. ']],38,54,0,71,0,8,263,0.08837209302325581,0.12558139534883722,0.16511627906976745,0.002325581395348837,0.0,0.21627906976744185,1,"['www.ons.gov', 'www.metoffice.gov', 'www.gov', 'www.statistics.gov', 'legislation.gov', 'www.ons.gov', 'wales.gov', 'statswales.gov', 'coflein.gov', 'www.number10.gov', 'www.gov', 'webarchive.nationalarchives.gov', 'wales.gov', 'www.royalmint.gov', 'www.statistics.gov', 'www.legislation.gov', 'www.gov', 'statswales.gov', 'www.justice.gov', 'www.ons.gov', '(www.statistics.gov', 'new.wales.gov', 'www.statswales.wales.gov', 'www.ons.gov', 'coflein.gov', 'www.ons.gov', 'www.ons.gov', 'wales.gov', 'wales.gov', 'new.wales.gov', 'morgangriffith.house.gov', 'wales.gov', 'nla.gov', 'wales.gov', 'law.gov', 'www.wales.gov', 'www.metoffice.gov', 'www.ons.gov', 'statswales.gov', 'new.wales.gov', 'wales.gov', 'www.legislation.gov', 'www.hmcourts-service.gov', 'webarchive.nationalarchives.gov', 'wales.gov', 'webarchive.nationalarchives.gov', 'www.metoffice.gov', 'www.statswales.wales.gov', 'statistics.gov', 'www.ons.gov', 'wales.gov', 'legislation.gov', 'webarchive.nationalarchives.gov', 'www.ons.gov', 'books.google.com', 'www.glamorgancricket.com', 'books.google.com', 'hansard.millbanksystems.com', 'hansard.millbanksystems.com', 'www.itv.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.bbc.com', 'books.google.com', 'www.uefa.com', 'applewarrior.com', 'www.historic-uk.com', 'corporate.dwrcymru.com', 'books.google.com', 'newcriterion.com', 'books.google.com', 'www.visitwales.com', 'books.google.com', 'stateofwales.com', 'www.loudersound.com', 'canugwerin.com', 'afi.com', 'www.royalmint.com', 'books.google.com', 'books.google.com', 'www.wales.com', 'www.wales.com', 'www.halcrow.com', 'books.google.com', 'diversiton.com', 'www.corusgroup.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'www.welshpremier.com', 'www.cnn.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.epcrugby.com', '.com', 'snowdoniaguide.com', 'www.bing.com', 'books.google.com', 'books.google.com', 'www.timet.com', 'www.itv.com', 'books.google.com', 'books.google.com', 'thecgf.com', '.com', 'news.nationalgeographic.com', 'www.historic-uk.com', 'www.oxfordreference.com', 'www.classicfm.com', 'books.google.com', 'books.google.com', 'www.bbc.com', '.com', 'www.socialistunity.com', 'www.itv.com', 'www.bbcgoodfood.com', 'books.google.com', 'www.royalmint.com', 'books.google.com', 'www.cardiff-airport.com', 'wales.com', 'www.shropshirestar.com', 'www.bbc.com', 'fraserofallander.org', 'hdi.globaldatalab.org', 'whc.unesco.org', 'www.iiss.org', 'www.ggat.org', 'www.iso.org', 'assemblywales.org', 'wayback.archive-it.org', 'www.byig-wlb.org', 'www.archiveswales.org', 'www.instituteforgovernment.org', 'www.rspb.org', 'www.agor.org', 'www.cartography.org', 'www.assemblywales.org', 'www.archiveswales.org', 'www.webarchive.org', 'www.rspb.org', 'www.sportwales.org', 'rspb.org', 'www.assemblywales.org', 'www.gweini.org', 'roads.org', 'llgc.org', 'newadvent.org', 'www.wbti.org', 'runeberg.org', 'www.ggat.org', 'www.planetmagazine.org', 'www.cllc.org', 'www.rcaconwy.org', 'www.llgc.org', 'assemblywales.org', 'gtj.org', 'www.webarchive.org', 'stamfordhistory.org', 'www.ggat.org', 'www.ggat.org', ['q. j. geol. soc. lond. ']]",69894,Require autoconfirmed or confirmed access (no expiry set),226867,1 September 2001,Asa~enwiki ,10608,129,2001-09-01,2001-09,2001
149,149,Lhoba people,https://en.wikipedia.org/wiki/Lhoba_people,19,0,"[None, None, None, None, None, None, None, None, None]","[['university of california at berkeley '], ['rajiv gandhi university via shodhganga '], ['jawaharlal nehru college']]",1,1,0,5,0,0,9,0.05263157894736842,0.05263157894736842,0.2631578947368421,0.0,0.0,0.10526315789473684,3,"['in.gov', 'books.google.com', 'books.google.com', 'www.indiandefencereview.com', 'www.north-east-india.com', 'www.dailypioneer.com', 'en.chinaculture.org', ['university of california at berkeley '], ['rajiv gandhi university via shodhganga '], ['jawaharlal nehru college']]",153035,Allow all users (no expiry set),18369,29 November 2002,Danny ,352,2,2002-11-29,2002-11,2002
150,150,Andhra Pradesh,https://en.wikipedia.org/wiki/Andhra_Pradesh,232,1,"['10.1017/s0026749x00004996', None, None]",[['[[modern asian studies']],13,43,0,111,0,0,66,0.05603448275862069,0.1853448275862069,0.47844827586206895,0.004310344827586207,0.0,0.24568965517241378,1,"['www.ap.gov', 'www.narl.gov', 'www.ap.gov', 'ap.gov', 'www.aponline.gov', 'www.censusindia.gov', 'www.ap.gov', 'aponline.gov', 'apedb.gov', 'www.censusindia.gov', 'www.ndrdgh.gov', 'dopr.gov', 'www.aponline.gov', 'www.censusindia.gov', 'nationalmap.gov', 'www.ap.gov', 'www.apgenco.gov', 'www.ap.gov', 'pib.gov', 'bse.ap.gov', 'www.aptransco.gov', 'www.ap.gov', 'www.aponline.gov', 'apsrtc.gov', 'bieap.gov', 'www.ap.gov', 'ap.gov', 'censusindia.gov', 'www.indianrailways.gov', 'www.aptdc.gov', 'www.ap.gov', 'www.caa.gov', 'www.ap.gov', 'www.scr.indianrailways.gov', 'www.ap.gov', 'aponline.gov', 'www.indiabudget.gov', 'www.ap.gov', 'ap.gov', 'www.portal.gsi.gov', 'studentinfo.ap.gov', 'schooledu.ap.gov', 'www.ap.gov', 'preethika.wordpress.com', 'guinnessworldrecords.com', 'timesofindia.indiatimes.com', 'deccan-journal.com', 'quickgs.com', 'books.google.com', 'www.newindianexpress.com', 'books.google.com', 'www.thehindu.com', 'www.newindianexpress.com', 'mapsofindia.com', 'www.thehindu.com', 'www.thehindubusinessline.com', 'zeenews.india.com', 'www.thehindu.com', 'www.thehindubusinessline.com', 'www.thehindu.com', 'www.thehindu.com', 'amaravativoice.com', 'www.thehindubusinessline.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.britannica.com', 'books.google.com', 'm.timesofindia.com', 'statisticstimes.com', 'www.newindianexpress.com', 'www.britannica.com', 'timesofindia.indiatimes.com', 'www.ndtv.com', 'www.asiantribune.com', 'www.thehindu.com', 'indiascanner.com', 'cleantechnica.com', 'deccanchronicle.com', 'www.populationu.com', 'www.sakshi.com', 'www.britannica.com', 'www.thehindu.com', 'www.travelandleisure.com', 'www.mid-day.com', 'www.britannica.com', 'books.google.com', 'gangavaram.com', 'books.google.com', 'www.thehindu.com', 'www.deccanchronicle.com', 'www.thehindu.com', 'www.thehindubusinessline.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'www.time.com', 'www.ndtv.com', 'news.google.com', 'www.forbes.com', 'www.thehindu.com', 'www.newindianexpress.com', 'books.google.com', 'www.deccanchronicle.com', 'books.google.com', 'www.thenewsminute.com', 'www.business-standard.com', 'www.thehindu.com', 'mihira.com', 'books.google.com', 'books.google.com', 'www.deccanchronicle.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehansindia.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.newindianexpress.com', 'www.thehindu.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.thehindubusinessline.com', 'books.google.com', 'english.sakshi.com', 'www.apassemblylive.com', 'www.indiatvnews.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'inc42.com', 'ndtv.com', 'books.google.com', 'www.tourisminap.com', 'www.andhraports.com', 'jagranjosh.com', 'ndtv.com', 'www.newindianexpress.com', 'andhrapradesh.pscnotes.com', 'www.templenet.com', 'deccanchronicle.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'www.ndtv.com', 'deccanchronicle.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'www.vizagport.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.nio.org', 'hdi.globaldatalab.org', 'www.isro.org', 'www.apsche.org', 'www.ramsar.org', 'www.rbi.org', 'isro.org', 'bseap.org', 'www.aplegislature.org', 'www.ctri.org', 'www.dghindia.org', 'ccrhindia.org', 'bseap.org', ['[[modern asian studies']]",2377,Allow all users (no expiry set),154169,29 October 2001,Tsja ,13822,63,2001-10-29,2001-10,2001
151,151,Serbia,https://en.wikipedia.org/wiki/Serbia,458,15,"['10.2298/gei1701127t', '10.1371/journal.pbio.2004956', '10.1080/21599165.2018.1490272', '10.1353/ser.2011.0038', '10.1016/j.jhevol.2011.03.003', '10.2298/eka1403029r', '10.4000/balkanologie.774', '10.1038/s41467-020-19493-3', '10.1080/1070289x.2014.969269', '10.17651/polon.37.9', '10.4467/25444654spp.19.004.10147', '10.1080/23745118.2017.1419599', '10.2298/vsp120205002s', '10.1080/13510347.2020.1758670', '10.3998/mp.9460447.0002.203', None, '29672508', None, None, '21507461', None, None, '33293507', None, None, None, None, '25536810', None, None, None, '5908072', None, None, None, None, None, '7723057', None, None, None, None, None, None, None]","[['glasnik etnografskog instituta sanu'], ['plos biology'], ['east european politics'], ['serbian studies'], ['journal of human evolution '], ['economic annals'], ['balkanologie. revue d'], ['nature communications'], [' identities'], ['polonica '], ['studia z zakresu prawa pracy i polityki społecznej'], ['european politics and society '], ['vojnosanit pregl '], ['democratization '], ['music and politics']]",45,56,0,163,0,1,179,0.0982532751091703,0.1222707423580786,0.3558951965065502,0.03275109170305677,0.0,0.25327510917030566,15,"['publikacije.stat.gov', 'www.siepa.gov', 'www.cia.gov', 'srbija.gov', 'www.mod.gov', 'www.export.gov', 'www.ekonomskitim.sr.gov', 'www.hidmet.gov', 'www.cia.gov', 'www.parlament.gov', 'www.mfa.gov', 'siepa.gov', 'www.mfa.gov', 'stat.gov', 'cia.gov', 'publikacije.stat.gov', 'www.loc.gov', 'parlament.gov', 'pod2.stat.gov', 'siepa.gov', 'www.stat.gov', 'www.trade.gov', 'www.mfa.gov', 'publikacije.stat.gov', 'mod.gov', 'www.mfa.gov', 'earthobservatory.nasa.gov', 'www.cia.gov', 'publikacije.stat.gov', 'pod2.stat.gov', 'siepa.gov', 'belgrade.usembassy.gov', 'stat.gov', 'publikacije.stat.gov', 'publikacije.stat.gov', 'www.arhivyu.gov', 'www.mfa.gov', 'siepa.gov', 'www.srbija.gov', 'www.cia.gov', 'www.srbija.gov', 'pod2.stat.gov', 'www.economy.gov', 'pod2.stat.gov', 'www.javnidug.gov', 'www.rik.parlament.gov', 'webrzs.stat.gov', 'www.srbija.gov', 'www.cia.gov', 'www.hidmet.gov', 'pod2.stat.gov', 'stat.gov', 'srbija.gov', 'bia.gov', 'siepa.gov', 'www.srbija.gov', 'books.google.com', 'books.google.com', 'www.serbianmonitor.com', 'books.google.com', 'rs.n1info.com', 'books.google.com', 'www.zumberacki-vikarijat.com', 'www.pfistudios.com', 'firstworldwar.com', 'books.google.com', 'www.nytimes.com', 'www.vreme.com', 'liberalniforum.com', 'books.google.com', 'sports.espn.go.com', 'balkans360.com', 'www.ft.com', 'books.google.com', 'today.in-24.com', 'www.carlsberggroup.com', 'www.exyuaviation.com', 'www.bbc.com', 'books.google.com', 'www.turorama.com', 'www.bbc.com', 'www.hartford-hwp.com', 'www.thebalkansdaily.com', 'uk.practicallaw.com', 'www.bbc.com', 'news.yahoo.com', 'www.xinhuanet.com', 'books.google.com', 'worldpopulationreview.com', 'books.google.com', 'www.pregled-rs.com', 'books.google.com', 'timesmachine.nytimes.com', 'amsglossary.allenpress.com', 'balkaninsight.com', 'intellinews.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.worldriskreport.com', 'books.google.com', 'books.google.com', 'www.cnn.com', 'books.google.com', 'books.google.com', 'bturn.com', 'www.aljazeera.com', 'rs.n1info.com', 'rs.n1info.com', 'books.google.com', 'medium.com', 'www.serbia-visit.com', 'balkaninsight.com', 'bitef.com', 'books.google.com', 'seenews.com', 'www.serbianrailways.com', 'balkaninsight.com', 'www.brewer-world.com', 'rs.n1info.com', 'books.google.com', 'books.google.com', 'rs.n1info.com', 'britannica.com', 'books.google.com', 'www.serbianmonitor.com', 'books.google.com', 'ogj.com', 'www.football-observatory.com', 'khazars.com', 'worldatlas.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.serbianmonitor.com', 'www.bbc.com', 'www.nysun.com', '2fwww.sacred-fr.com', 'seenews.com', 'books.google.com', 'books.google.com', 'euobserver.com', 'books.google.com', 'books.google.com', 'rs.n1info.com', 'books.google.com', 'books.google.com', 'au.totaltravel.yahoo.com', 'belgraded.com', 'abcnews.go.com', 'ww1live.wordpress.com', 'www.bastabalkana.com', 'wrmjournal.com', 'timesofindia.indiatimes.com', 'soccerlens.com', 'muzejirade.com', 'www.google.com', 'books.google.com', 'www.kosovopolice.com', 'books.google.com', 'www.britannica.com', 'www.reuters.com', 'serbia.com', 'books.google.com', 'www.pregled-rs.com', 'books.google.com', 'pqasb.pqarchiver.com', 'bturn.com', 'www.vesti-online.com', 'www.earthsendangered.com', 'turistickimagazin.com', 'www.ekapija.com', 'kustu.com', 'rememberingyugoslavia.com', 'books.google.com', 'books.google.com', 'joakimvujic.com', 'myforevertravel.com', 'rs.n1info.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.alexa.com', 'rs.n1info.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'www.srbijagas.com', 'www.dipublico.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.beogradskisajamknjiga.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.huffingtonpost.com', 'books.google.com', 'www.bulgaria-italia.com', 'www.ch-aviation.com', 'www.britannica.com', 'www.shanghairanking.com', 'books.google.com', 'serbia-times.com', 'filmneweurope.com', 'knoema.com', 'books.google.com', 'theculturetrip.com', 'danube-cooperation.com', 'books.google.com', 'rs.n1info.com', 'balkangreenenergynews.com', 'books.google.com', 'www.calvertjournal.com', 'rs.n1info.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.sgd.org', 'yadvashem.org', 'discoverserbia.org', 'www.kinoteka.org', 'www.batut.org', 'www.unesco.org', 'www.imf.org', 'www.kinoteka.org', 'www.fifoost.org', 'openknowledge.worldbank.org', 'www.socialprogress.org', 'iucn.org', 'uvac.org', 'collection.cooperhewitt.org', 'www.worldenergy.org', 'seecult.org', 'www.globalsecurity.org', 'imf.org', 'www.exitfest.org', 'waterpoloserbia.org', 'web.worldbank.org', 'rsf.org', 'faostat3.fao.org', 'hdr.undp.org', 'www.osce.org', 'www.visitserbia.org', 'imf.org', 'www.amnesty.org', 'www.freedomhouse.org', 'humanrightshouse.org', 'www.ccre.org', 'zeno.org', 'www.pbs.org', 'www.rra.org', 'ei-ie.org', 'www.visionofhumanity.org', 'wayback.archive-it.org', 'ourworldindata.org', 'www.turizamprijepolje.org', 'exitfest.org', 'www.rferl.org', 'combatgenocide.org', 'www.slobodnaevropa.org', 'www.worldbank.org', 'royalfamily.org', ['glasnik etnografskog instituta sanu'], ['plos biology'], ['east european politics'], ['serbian studies'], ['journal of human evolution '], ['economic annals'], ['balkanologie. revue d'], ['nature communications'], [' identities'], ['polonica '], ['studia z zakresu prawa pracy i polityki społecznej'], ['european politics and society '], ['vojnosanit pregl '], ['democratization '], ['music and politics']]",29265,Require administrator access (no expiry set),272426,15 December 2001,David Parker ,17030,35,2001-12-15,2001-12,2001
152,152,Scotland,https://en.wikipedia.org/wiki/Scotland,423,5,"['10.1127/zfg/30/1987/407', '10.1093/acref/9780199545568.001.0001', '10.1215/00982601-29-2-25', '10.1080/713999852', None, None, None, None, None, None, None, None]","[['[[zeitschrift für geomorphologie'], ['oxford university press'], ['eighteenth-century life '], ['culture']]",39,85,0,63,0,7,224,0.09219858156028368,0.20094562647754138,0.14893617021276595,0.01182033096926714,0.0,0.3049645390070922,4,"['www.ons.gov', 'www.opsi.gov', 'www.scotcourts.gov', 'www.gov', 'www.gov', 'www.gov', 'www.legislation.gov', 'www.legislation.gov', 'www.scotlandscensus.gov', 'scot.gov', 'nitakeacloserlook.gov', 'www.opsi.gov', 'www.metoffice.gov', 'www.scotlandscensus.gov', 'www.gov', 'www.gov', 'www.nrscotland.gov', 'firstminister.gov', 'www.metoffice.gov', 'www.gov', 'www.gov', 'www.ons.gov', 'www.gov', 'www.gov', 'www.nationalarchives.gov', 'ons.gov', 'www.gov', 'dataportal.orr.gov', 'www.metoffice.gov', 'www.gov', 'www.scotlandscensus.gov', 'www.scotlandoffice.gov', 'www.gov', 'www.saas.gov', 'cosla.gov', 'www.gov', 'www.gov', 'beta.gov', 'www.gov', 'www.gov', 'www.gov', 'www.gov', 'www.gov', 'dca.gov', 'beta.gov', 'beta.gov', 'www.forestry.gov', 'nationalarchives.gov', 'www.gov', 'www.scotland.gov', 'www.ons.gov', 'www.gov', 'cosla.gov', 'www.opsi.gov', 'www.gov', 'www.nationalarchives.gov', 'www.gov', 'www.gov', 'www.ons.gov', 'www.rail-reg.gov', 'transport.gov', 'www.gov', 'factfinder.census.gov', 'sps.gov', 'www.gov', 'www.number10.gov', 'www.transport.gov', 'cosla.gov', 'www.gov', 'www.nas.gov', 'www.gov', 'www.nas.gov', 'www.scotlandscensus.gov', 'www.gov', 'scotland.gov', 'www.gov', 'www.nrscotland.gov', 'scotlandscensus.gov', 'factfinder.census.gov', 'www.scotlandscensus.gov', 'www.nationalarchives.gov', 'www.legislation.gov', 'www.scotlandscensus.gov', 'dca.gov', 'www.gov', 'www.pgatour.com', 'www.festival-interceltique.com', 'www.historyscotland.com', 'books.google.com', '90min.com', 'www.bbc.com', 'www.timeshighereducation.com', 'www.britannica.com', 'rampantscotland.com', 'www.bbcstudios.com', 'scotsman.com', 'www.bbc.com', 'books.google.com', 'news.scotsman.com', 'news.google.com', 'heraldscotland.com', 'www.celticconnections.com', 'books.google.com', 'www.bbc.com', 'breakingnews.heraldscotland.com', 'books.google.com', 'americanheritage.com', 'www.pgatour.com', 'news.scotsman.com', 'www.britannica.com', 'fifa.com', 'rampantscotland.com', 'intheknowtraveler.com', 'www.scottishlegal.com', 'www.scotsman.com', 'www.itv.com', 'thestudiomap.com', 'books.google.com', 'www.historichighlanders.com', 'newtonmore.com', 'www.newstatesman.com', 'espn.com', 'www.newsnetscotland.com', 'books.google.com', 'www.fifa.com', 'scotsman.com', 'www.scotsman.com', 'www.heraldscotland.com', 'www.scotsman.com', 'bbc.com', 'powells.com', 'www.historic-uk.com', 'ca.encarta.msn.com', 'www.holyrood.com', 'time.com', 'visitscotland.com', 'books.google.com', 'www.bbc.com', 'fifa.com', 'www.heraldscotland.com', 'scottishfinancialreview.com', 'www.bbc.com', 'www.nationalcelticfestival.com', 'scottishhistorysociety.com', 'www.scotsman.com', 'www.taste-of-scotland.com', 'www.bbc.com', 'books.google.com', 'hdi.globaldatalab.org', 'www.scottishgolfhistory.org', 'www.historyofparliamentonline.org', 'scotland.org', 'www.catholic.org', 'www.treefestscotland.org', 'www.instituteforgovernment.org', 'rbge.org', 'www.lawscot.org', 'www.flaginstitute.org', 'www.britishirishcouncil.org', 'www.scotland.org', 'www.catholic.org', 'www.catholic.org', 'churchofscotland.org', 'churchofscotland.org', 'www.ltscotland.org', 'www.scan.org', 'www.lawscot.org', 'www.iso.org', 'www.britishirish.org', 'cgcs.org', 'www.catholic.org', 'snh.org', 'cgcs.org', 'assets.cambridge.org', 'archive.ifla.org', 'www.scis.org', 'www.carnegie-trust.org', 'www.scotland.org', 'www.scotch-whisky.org', 'www.scotland.org', 'www.rspb.org', 'scotland.org', 'www.scottishaffairs.org', 'www.scotland-malawipartnership.org', 'www.scotland.org', 'www.ltscotland.org', 'www.scotch-whisky.org', ['[[zeitschrift für geomorphologie'], ['oxford university press'], ['eighteenth-century life '], ['culture']]",26994,Require administrator access (no expiry set),236235,1 October 2001,Clasqm ,17332,33,2001-10-01,2001-10,2001
153,153,United Kingdom,https://en.wikipedia.org/wiki/United_Kingdom,684,24,"['10.1080/0031322x.1996.9970192', '10.1080/01419870701599465', '10.1177/0038038511419195', '10.1093/publius/pjj011', '10.1093/oxfordjournals.pubjof.a029948', '10.1086/644536', '10.1038/s41467-020-19493-3', '10.1093/pa/52.1.19', '10.1098/rspb.2006.3627', 'abs/10.1080/04597222.2021.1868791?journalcode=tmib20', '10.1111/1468-2230.00203', '10.1098/rspa.1948.0129', '10.1080/21622671.2021.1921613', '10.1177/20419058211000996', '10.1093/slr/hmab003/6213886', '10.1093/icon/2.3.545', '10.1038/159297a0', '10.1080/13501763.2021.1876156', '10.1093/biosci/bix014', None, None, None, None, None, None, '33293507', None, '17002951', None, None, None, None, None, None, None, None, None, '28608869', None, None, None, None, None, None, '7723057', None, '1635457', None, None, None, None, None, None, None, None, None, '5451287']","[['patterns of prejudice'], ['ethnic and racial studies'], ['sociology'], ['publius'], ['publius'], ['journal of british studies'], ['nature communications'], ['parliamentary affairs'], ['proceedings of the royal society b'], [' the military balance'], ['the modern law review'], ['proceedings of the royal society of london'], ['territory', '[[taylor '], ['[[sage publishing', 'political insight '], ['[[statute law review', '[[oxford university press'], ['international journal of constitutional law'], ['nature'], ['[[journal of european public policy', '[[taylor '], ['bioscience']]",67,113,0,166,0,15,299,0.097953216374269,0.1652046783625731,0.24269005847953215,0.03508771929824561,0.0,0.2982456140350877,19,"['www.statistics.gov', 'www.cia.gov', 'history.blog.gov', 'archive.defra.gov', 'www.gov', 'www.ons.gov', 'www.dft.gov', 'www.gov', 'webarchive.nationalarchives.gov', 'www.royal.gov', 'www.ons.gov', 'www.statistics.gov', 'www.ons.gov', 'www.cia.gov', 'webarchive.nationalarchives.gov', 'www.northernireland.gov', 'www.bis.gov', 'webarchive.nationalarchives.gov', 'www.statistics.gov', 'webarchive.nationalarchives.gov', 'www.ons.gov', 'www.ons.gov', 'webarchive.nationalarchives.gov', 'webarchive.nationalarchives.gov', 'www.gov', 'www.gov', 'www.ons.gov', 'www.ukba.homeoffice.gov', 'www.gov', 'www.gov', 'www.scotcourts.gov', 'ukclimateprojections.metoffice.gov', 'ons.gov', 'www.gos.gov', 'www.ons.gov', 'assets.publishing.service.gov', 'orr.gov', 'www.scotlandscensus.gov', 'www.scotcourts.gov', 'www.nationalarchives.gov', 'www.culture.gov', 'www.lga.gov', 'www.gov', 'ons.gov', 'www.ons.gov', 'www.ons.gov', 'www.northernireland.gov', 'www.gov', 'assets.publishing.service.gov', 'www.ons.gov', 'www.statistics.gov', 'webarchive.nationalarchives.gov', 'www.cia.gov', 'www.justice.gov', 'www.ons.gov', 'www.ons.gov', 'assets.publishing.service.gov', 'www.environment-agency.gov', 'www.eia.gov', 'www.statistics.gov', 'www.royalinsight.gov', 'www.ons.gov', 'webarchive.nationalarchives.gov', 'tonto.eia.doe.gov', 'www.gov', 'www.gov', 'www.nationalarchives.gov', 'webarchive.nationalarchives.gov', 'www.eia.gov', 'www.gov', 'www.royal.gov', 'www.statistics.gov', 'orr.gov', 'www.statistics.gov', 'www.ons.gov', 'www.statistics.gov', 'www.gov', 'www.gov', 'obamawhitehouse.archives.gov', 'www.eia.gov', 'www.gro-scotland.gov', 'neighbourhood.statistics.gov', 'www.london.gov', 'www.ons.gov', 'www.gov', 'www.ons.gov', 'www.cia.gov', 'www.ons.gov', 'www.ons.gov', 'college-of-arms.gov', 'www.direct.gov', 'www.cia.gov', 'www.cia.gov', 'webarchive.nationalarchives.gov', 'www.eia.gov', 'www.gov', 'www.coal.gov', 'www.scotcourts.gov', 'www.ons.gov', 'www.gov', 'www.gov', 'www.gov', 'www.culture.gov', 'www.ons.gov', 'www.gov', 'www.loc.gov', 'www.gov', 'www.neighbourhood.statistics.gov', 'www.ons.gov', 'www.census.gov', 'webarchive.nationalarchives.gov', 'www.gov', 'assets.publishing.service.gov', 'www.britannica.com', 'books.google.com', 'traveltips.usatoday.com', 'www.topuniversities.com', 'railway-technology.com', 'www.ukmediacentre.pwc.com', 'books.google.com', 'www.washingtonpost.com', 'books.google.com', 'deutschebahn.com', 'www.trevorharley.com', 'www.forbes.com', 'www.bbc.com', 'www.nytimes.com', 'en.oxforddictionaries.com', 'www.ft.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'www.oxfordreference.com', 'www.bcg.com', 'edition.cnn.com', 'books.google.com', 'www.forbes.com', 'learnersdictionary.com', 'www.llrx.com', 'www.rlwc08.com', 'www.oxfordmusiconline.com', 'books.google.com', 'www.zyen.com', 'books.google.com', 'equalityhumanrights.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'indexmundi.com', 'www.bbc.com', 'books.google.com', 'atlapedia.com', 'uk.reuters.com', 'books.google.com', 'www.stockmarketwire.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.reuters.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.time.com', 'books.google.com', 'www.fifa.com', 'www.medianewsline.com', 'www.timeshighereducation.com', 'allmusic.com', 'news.scotsman.com', 'books.google.com', 'www.statista.com', 'books.google.com', 'newsfeed.time.com', 'www.playbillarts.com', 'books.google.com', 'www.eurotunnel.com', 'www.google.com', 'books.google.com', 'www.com', 'rollingstone.com', 'books.google.com', 'www.shanghairanking.com', 'edition.cnn.com', 'www.britannica.com', 'www.oxforddictionaries.com', 'encyclopedia2.thefreedictionary.com', 'www.internetworldstats.com', 'cibc.com', 'uk.practicallaw.thomsonreuters.com', 'www.emimusic.com', 'www.medianewsline.com', 'books.google.com', 'www.allmusic.com', 'books.google.com', 'www.statista.com', 'bbc.com', 'books.google.com', 'itv.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.economist.com', 'books.google.com', 'books.google.com', 'www.emimusic.com', 'www.bbc.com', 'www.bloomberg.com', 'www.bbc.com', 'news.nationalgeographic.com', 'www.euromonitor.com', 'www.ealingstudios.com', 'books.google.com', 'books.google.com', 'niwater.com', 'www.statista.com', 'books.google.com', 'books.google.com', 'encarta.msn.com', 'globescan.com', 'books.google.com', 'books.google.com', 'www.wales.com', 'books.google.com', 'www.britannica.com', 'www.pgatour.com', 'books.google.com', 'www.trevorharley.com', 'books.google.com', 'www.equalityhumanrights.com', 'www.theaustralian.com', 'www.itftennis.com', 'books.google.com', 'books.google.com', 'www.allmusic.com', 'www.scotsman.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.newscorp.com', 'www.newscorp.com', 'www.ipsos-mori.com', 'books.google.com', 'www.redbull.com', 'books.google.com', 'books.google.com', 'www.billboard.com', 'books.google.com', 'www.encyclopedia.com', 'www.ft.com', 'www.nme.com', 'www.allmusic.com', 'www.usnews.com', 'www.cnn.com', 'books.google.com', 'finance.yahoo.com', 'encarta.msn.com', 'books.google.com', 'www.mastercard.com', 'www.britannica.com', 'www.oxfordmusiconline.com', 'books.google.com', 'www.migrationwatchuk.com', 'books.google.com', 'www.bbc.com', 'bbc.com', 'www.billboard.com', 'www.collinsdictionary.com', 'books.google.com', 'www.redorbit.com', 'books.google.com', 'www.instituteforgovernment.org', 'unstats.un.org', 'www.oecd.org', 'www.wssinfo.org', 'www.britishcouncil.org', 'www.churchofscotland.org', 'stakeholders.ofcom.org', 'www.ltscotland.org', 'www.healthp.org', 'news.adventist.org', 'www.migrationwatchuk.org', 'royalsociety.org', 'www.npr.org', 'www.ccea.org', 'www.sqa.org', 'www.scis.org', 'unstats.un.org', 'olympic.org', 'ourworldindata.org', 'nobelprize.org', 'data.imf.org', 'www.thecommonwealth.org', 'www.ukotcf.org', 'www.iso.org', 'runeberg.org', 'www.migrationinformation.org', 'www.gmb.org', 'www.scotland.org', 'www.ippr.org', 'www.cartography.org', 'internationaltransportforum.org', 'www.chathamhouse.org', 'us.oecd.org', 'www.imf.org', 'scotland.org', 'www.mersey-gateway.org', 'www.foe-scotland.org', 'hdr.undp.org', 'www.tate.org', 'esa.un.org', 'www.imf.org', 'www.thecommonwealth.org', 'www.world-nuclear.org', 'www.unesco.org', 'www.commonwealthofnations.org', 'www.sipri.org', 'dictionary.cambridge.org', 'www.wssinfo.org', 'www.world-tourism.org', 'www.bfi.org', 'www.instituteforgovernment.org', 'portal.unesco.org', 'www.prisonstudies.org', 'www.cofe.anglican.org', 'databank.worldbank.org', 'www.seaaroundus.org', 'data.un.org', 'www.ofcom.org', 'www.literaturewales.org', 'www.royal-navy.org', 'www.scotland.org', 'archontology.org', 'rooseveltinstitute.org', 'www.ukfilmcouncil.org', 'commons.wikimedia.org', 'stats.oecd.org', 'www.internationalpublishers.org', ['patterns of prejudice'], ['ethnic and racial studies'], ['sociology'], ['publius'], ['publius'], ['journal of british studies'], ['nature communications'], ['parliamentary affairs'], ['proceedings of the royal society b'], [' the military balance'], ['the modern law review'], ['proceedings of the royal society of london'], ['territory', '[[taylor '], ['[[sage publishing', 'political insight '], ['[[statute law review', '[[oxford university press'], ['international journal of constitutional law'], ['nature'], ['[[journal of european public policy', '[[taylor '], ['bioscience']]",31717,Require administrator access (no expiry set),353061,2 November 2001,195.70.85.xxx ,25230,67,2001-11-02,2001-11,2001
154,154,Hungary,https://en.wikipedia.org/wiki/Hungary,269,7,"['10.1080/13510347.2021.1922390', '10.1093/biosci/bix014', '10.1017/s0020818300035414', '10.1038/s41467-020-19493-3', '10.1787/data-00544-en', None, '28608869', None, '33293507', None, None, '5451287', None, '7723057', None]","[['democratization '], ['bioscience'], ['international organization'], ['nature communications'], ['oecd health statistics ']]",25,14,0,77,0,3,145,0.09293680297397769,0.05204460966542751,0.2862453531598513,0.026022304832713755,0.0,0.17100371747211895,5,"['www.cia.gov', 'www.mfa.gov', 'www.cia.gov', 'nkfih.gov', 'lcweb2.loc.gov', 'www.cia.gov', 'www.cia.gov', 'cia.gov', 'www.cia.gov', 'www.cia.gov', 'lcweb2.loc.gov', 'www.mfa.gov', 'www.cia.gov', 'www.cia.gov', 'www.startupranking.com', 'books.google.com', 'hungarianhistory.com', 'www.euronews.com', 'www.economistinsights.com', 'fifa.com', 'books.google.com', 'imtj.com', 'books.google.com', 'www.bbc.com', 'geography.about.com', 'books.google.com', 'books.google.com', 'www.digitaljournal.com', 'ratings.fide.com', 'www.britannica.com', 'www.hungarianhistory.com', 'books.google.com', 'soccernet.espn.go.com', 'ukmediacentre.pwc.com', 'hungarianfreepress.com', 'books.google.com', 'www.fia.com', 'www.forbes.com', 'books.google.com', 'books.google.com', 'geocities.com', 'books.google.com', 'asiatravel.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'medalspercapita.com', 'www.gptoday.com', 'soccernet.espn.go.com', 'books.google.com', 'www.encyclopedia.com', 'www.cnbc.com', 'hungarianhistory.com', 'money.cnn.com', 'findarticles.com', 'historicaltextarchive.com', 'books.google.com', 'books.google.com', 'www.fifa.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.as.com', 'budapestcorner.com', 'books.google.com', 'books.google.com', 'imtj.com', 'books.google.com', 'books.google.com', 'books.google.com', 'dw.com', 'www.bbc.com', 'www.time.com', 'medalspercapita.com', 'budapestagent.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.tamupress.com', 'www.bloomberg.com', 'www.ft.com', 'hngary.com', 'query.nytimes.com', 'www.britannica.com', 'britannica.com', 'www.royal-tokaji.com', 'stats.oecd.org', 'hdr.undp.org', 'www.globalinnovationindex.org', 'magyarnews.org', 'www.jdc.org', 'visionofhumanity.org', 'fao.org', 'www3.weforum.org', 'www.globalinnovationindex.org', 'www.ushmm.org', 'freedomhouse.org', 'www.npr.org', 'climate-data.org', 'ourworldindata.org', 'www.constituteproject.org', 'ushmm.org', 'www.unevoc.unesco.org', 'portal.unesco.org', 'www.imf.org', 'www.jstor.org', 'web.worldbank.org', 'data.worldbank.org', 'www.h-net.org', 'eliznik.org', 'www.imf.org', ['democratization '], ['bioscience'], ['international organization'], ['nature communications'], ['oecd health statistics ']]",13275,Allow all users (no expiry set),221062,9 May 2001,63.115.18.xxx ,13424,23,2001-05-09,2001-05,2001
155,155,Greece,https://en.wikipedia.org/wiki/Greece,382,11,"['10.1093/biosci/bix014', '10.1179/byz.1999.23.1.195', '10.1017/s0018246x00026200', '10.5070/c311008864', '10.12681/mnimon.171', '10.1080/14623520801950820', '10.1038/s41586-019-1376-z', '10.12681/mnimon.735', '10.4000/ceb.835', '10.1038/s41467-020-19493-3', '10.1080/01402380512331341121', '28608869', None, None, None, None, None, '31292546', None, None, '33293507', None, '5451287', None, None, None, None, None, None, None, None, '7723057', None]","[['bioscience'], ['byzantine and modern greek studies'], ['the historical journal'], ['california italian studies'], ['μνήμων'], [' journal of genocide research '], ['[[nature '], ['μνήμων'], ['cahiers balkaniques'], ['nature communications'], ['[[west european politics ']]",38,11,0,154,0,7,161,0.09947643979057591,0.028795811518324606,0.4031413612565445,0.028795811518324606,0.0,0.15706806282722513,11,"['www.cia.gov', '2009-2017.state.gov', 'www.cia.gov', 'rita.dot.gov', '2001-2009.state.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.investingreece.gov', 'cia.gov', 'www.cia.gov', 'culinarybackstreets.com', 'books.google.com', 'www.bloomberg.com', 'www.youtube.com', 'www.reuters.com', 'books.google.com', 'greeka.com', 'books.google.com', 'books.google.com', 'www.dw.com', 'books.google.com', 'www.fiba.com', 'books.google.com', 'www.economist.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.bloomberg.com', 'books.google.com', 'www.reuters.com', 'www.nytimes.com', 'www.ethnologue.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.openjourney.com', 'euobserver.com', 'www.euromoney.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'dw.com', 'www.euromoney.com', 'www.ekathimerini.com', 'books.google.com', 'www.ft.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.ekathimerini.com', 'www.fifa.com', 'culinarybackstreets.com', 'www.economist.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'books.google.com', 'www.aljazeera.com', 'www.highbeam.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.bloomberg.com', 'books.google.com', 'www.smithsonianmag.com', 'books.google.com', 'books.google.com', 'www.bbc.com', 'books.google.com', 'www.businessinsider.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'indexmundi.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'www.wsj.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.slate.com', 'books.google.com', 'books.google.com', 'sports.espn.go.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'www.newstatesman.com', 'books.google.com', 'www.ft.com', 'www.youtube.com', 'www.balkaninsight.com', 'books.google.com', 'books.google.com', 'www.bbc.com', 'www.bloomberg.com', 'www.reuters.com', 'www.ft.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', '24grammata.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'www.nytimes.com', 'books.google.com', 'www.bbc.com', 'books.google.com', 'www.britannica.com', 'www.lonelyplanet.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.reuters.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'www.bloomberg.com', 'egolpio.com', 'books.google.com', 'www.foreignaffairs.com', 'www.newsweek.com', 'www.ekathimerini.com', 'www.aljazeera.com', 'books.google.com', 'www.britannica.com', 'www.nytimes.com', 'books.google.com', 'www.bbc.com', 'www.travelandleisure.com', 'books.google.com', 'www.bbc.com', 'www.marketwatch.com', 'www.newsweek.com', 'www.usnews.com', 'www.qgazette.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'www.newsnowgr.com', 'www.travelandleisure.com', 'bruegel.org', 'download.jw.org', 'www.savethechildren.org', 'www.worldcat.org', 'data.worldbank.org', 'data.worldbank.org', 'stats.oecd.org', 'www.imf.org', 'wildhunt.org', 'www.pewforum.org', 'www.sbl-site.org', 'oecdbetterlifeindex.org', 'ourworldindata.org', 'w.oecdbetterlifeindex.org', 'data.worldbank.org', 'www.unwto.org', 'stats.oecd.org', 'www.migrationpolicy.org', 'www.wttc.org', 'whc.unesco.org', 'www.imf.org', 'www.imf.org', 'www.unctad.org', 'www.oecd.org', 'www.thisisathens.org', 'greece.org', 'data.unhcr.org', 'www.hri.org', 'www.unctad.org', 'hdr.undp.org', 'www.npr.org', 'data.worldbank.org', 'www.hri.org', 'hdr.undp.org', 'phys.org', 'www.unctad.org', 'www.imf.org', 'unstats.un.org', ['bioscience'], ['byzantine and modern greek studies'], ['the historical journal'], ['california italian studies'], ['μνήμων'], [' journal of genocide research '], ['[[nature '], ['μνήμων'], ['cahiers balkaniques'], ['nature communications'], ['[[west european politics ']]",12108,Require autoconfirmed or confirmed access (no expiry set),299993,10 September 2001,Koyaanis Qatsi ,19482,9,2001-09-10,2001-09,2001
156,156,Germany,https://en.wikipedia.org/wiki/Germany,290,16,"['10.1080/09668139408412190', '10.1038/nature07995', '10.1093/biosci/bix014', '10.2307/1498562', '10.1093/hwj/dbp009', '10.1093/ehr/ceq276', '10.1017/s0043887100002604', '10.1086/467481', '10.1073/pnas.1012722107', '10.1111/j.1468-229x.1934.tb01791.x', '10.2307/3113137', '10.1038/d41586-019-00910-7', '10.1177/002200949002500207', '10.1080/07075332.2005.9641060', '12288331', '19444215', '28608869', None, None, None, None, None, '21041630', None, None, '30918381', None, None, None, None, '5451287', None, None, None, None, None, '2993404', None, None, None, None, None]","[['europe-asia studies'], ['nature'], ['bioscience'], ['western folklore'], ['history workshop journal'], ['the english historical review'], ['world politics '], ['[[journal of legal studies'], ['[[proceedings of the national academy of sciences of the united states of america'], ['history '], ['the business history review '], ['nature'], ['journal of contemporary history'], ['the international history review']]",39,9,0,66,0,4,156,0.13448275862068965,0.03103448275862069,0.22758620689655173,0.05517241379310345,0.0,0.2206896551724138,14,"['germany.usembassy.gov', 'www.nationalarchives.gov', 'lcweb2.loc.gov', 'blogs.loc.gov', 'history.state.gov', 'www.eia.gov', 'www.archives.gov', 'www.cia.gov', 'www.state.gov', 'gizmodo.com', 'www.statista.com', 'www.statista.com', 'euractiv.com', 'www.nytimes.com', 'www.demographia.com', 'www.nytimes.com', 'www.statista.com', 'www.france24.com', 'www.devex.com', 'www.dw.com', 'www.bbc.com', 'www.bbc.com', 'airmundo.com', 'www.nytimes.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'theconversation.com', 'au.news.yahoo.com', 'www.ft.com', 'books.google.com', 'www.sciencealert.com', 'www.nytimes.com', 'www.dw.com', 'www.nytimes.com', 'www.nytimes.com', 'www.bbc.com', 'www.janes.com', 'www.dw.com', 'www.cnn.com', 'www.nasdaq.com', 'www.bloomberg.com', 'www.foodandwine.com', 'www.cnn.com', 'www.indexmundi.com', 'www.german-way.com', 'www.dw.com', 'thediplomat.com', 'www.statista.com', 'www.uefa.com', 'books.google.com', 'www.dw.com', 'books.google.com', 'www.topuniversities.com', 'www.timeshighereducation.com', 'www.fifa.com', 'www.electrive.com', 'www.statista.com', 'www.germanwineusa.com', 'www.dw.com', 'www.statista.com', 'www.fifa.com', 'www.britannica.com', 'm.timesofindia.com', 'www.dw.com', 'www.bbc.com', 'fortune.com', 'www.businessinsider.com', 'eurail.com', 'books.google.com', 'www.nytimes.com', 'www.dw.com', 'www.statista.com', 'www.theartnewspaper.com', 'www.imf.org', 'www.internationalpublishers.org', 'www.weforum.org', 'www.imf.org', 'germanlawarchive.iuscomp.org', 'www3.weforum.org', 'www.ushmm.org', 'internationalinsider.org', 'www.sipri.org', 'internationalinsider.org', 'www.cleanenergywire.org', 'data.oecd.org', 'www.ushmm.org', 'www.unesco.org', 'stats.oecd.org', 'www.wendemuseum.org', 'germanhistorydocs.ghi-dc.org', 'dataunodc.un.org', 'encyclopedia.ushmm.org', 'data.worldbank.org', 'wenr.wes.org', 'encyclopedia.ushmm.org', 'www.ambafrance-uk.org', 'medialandscapes.org', 'www.internationaltransportforum.org', 'www.un.org', 'germanfoods.org', 'www.cleanenergywire.org', 'hdr.undp.org', 'nobelprize.org', 'humanright2water.org', 'www.britishmuseum.org', 'www.sipri.org', 'www.transparency.org', 'whc.unesco.org', 'www.holocaustchronicle.org', 'www.holocaust-history.org', 'www.climateaction.org', 'data.worldbank.org', ['europe-asia studies'], ['nature'], ['bioscience'], ['western folklore'], ['history workshop journal'], ['the english historical review'], ['world politics '], ['[[journal of legal studies'], ['[[proceedings of the national academy of sciences of the united states of america'], ['history '], ['the business history review '], ['nature'], ['journal of contemporary history'], ['the international history review']]",11867,Require administrator access (no expiry set),197977,9 November 2001,Magnus Manske ,20372,30,2001-11-09,2001-11,2001
157,157,Abruzzo,https://en.wikipedia.org/wiki/Abruzzo,71,0,[],[],5,0,0,22,0,1,43,0.07042253521126761,0.0,0.30985915492957744,0.0,0.0,0.07042253521126761,0,"['www.resources.immobiliarecaserio.com', 'www.italyheritage.com', 'www.hotelposeidontortoreto.com', 'www.nytimes.com', 'www.liveandinvestoverseas.com', 'marinape.com', 'www.delallo.com', 'www.interamniaworldcup.com', 'www.lifeinabruzzo.com', 'en.com', 'www.abruzzoruralproperty.com', 'oliveoilsindia.com', 'books.google.com', 'www.academiabarilla.com', 'mariobatali.com', 'books.google.com', 'books.google.com', 'www.italy-schools.com', 'books.google.com', 'www.deliciousitaly.com', 'abruzzoairport.com', 'www.huffingtonpost.com', 'www.eib.org', 'hdi.globaldatalab.org', 'abruzzomoliseheritagesociety.org', 'www.eib.org', 'www.abruzzomoliseheritagesociety.org']",79460,Allow all users (no expiry set),72058,2 September 2002,64.59.222.4 ,1927,4,2002-09-02,2002-09,2002
158,158,France,https://en.wikipedia.org/wiki/France,530,7,"['10.2307/2610008', '10.1007/978-0-230-36688-6', '10.2105/ajph.2012.301136', '10.1038/s41467-020-19493-3', '10.1093/gao/9781884446054.article.t063666', '10.1016/j.trim.2007.03.002', 'pdf/10.18111/9789284421152', None, None, '23327250', '33293507', None, '17584595', None, None, None, '3673512', '7723057', None, None, None]","[['[[international affairs '], ['palgrave macmillan '], ['american journal of public health'], ['nature communications'], ['oxford university press'], ['transpl immunol. '], ['united nations world tourism organization ']]",93,11,0,181,0,8,230,0.17547169811320754,0.020754716981132074,0.34150943396226413,0.013207547169811321,0.0,0.20943396226415095,7,"['www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.nga.gov', 'www.cia.gov', '2001-2009.state.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'about.com', 'books.google.com', 'books.google.com', 'www.visualcapitalist.com', 'www.worldatlas.com', 'books.google.com', 'medoc-tourisme.com', 'h2g2.com', 'www.com', 'photius.com', 'www.scientificamerican.com', 'www.britannica.com', 'nakedtranslations.com', 'books.google.com', 'www.actu-environnement.com', 'www.statistiques-mondiales.com', 'www.france24.com', 'observatoire.ojd.com', 'www.3starrestaurants.com', 'www.reuters.com', 'books.google.com', 'nationmaster.com', 'books.google.com', 'www.usfunds.com', 'www.uefa.com', 'www.csmonitor.com', 'about-france.com', 'www.spglobal.com', 'about-france.com', 'www.globalpost.com', 'www.economist.com', 'www.forbes.com', 'www.laprovence.com', 'www.washingtonpost.com', 'www.globalgovernmentforum.com', 'www.nytimes.com', 'www.ojd.com', 'books.google.com', 'www.uciprotour.com', 'www.nytimes.com', 'whatsonwhen.com', 'www.usinenouvelle.com', 'books.google.com', 'www.nytimes.com', 'timeanddate.com', 'completelynovel.com', 'www.businessinsider.com', 'green.blogs.nytimes.com', 'www.frenchriviera-tourism.com', 'www.statista.com', 'www.britannica.com', 'www.britannica.com', 'www.secureworldexpo.com', 'afrik.com', 'www.natureindex.com', 'publications.credit-suisse.com', 'observatoire.ojd.com', 'europeupclose.com', 'www.irishtimes.com', 'www.intersurgtech.com', 'www.ey.com', 'www.123voyage.com', 'www.nytimes.com', 'www.bbc.com', 'myfrenchproperty.com', 'books.google.com', 'books.google.com', 'www.natureindex.com', 'books.google.com', 'www.themeit.com', 'www.britannica.com', 'www.ambest.com', 'www.scienceshumaines.com', 'www.britannica.com', 'www.nytimes.com', 'tourmag.com', 'intstudy.com', 'edition.cnn.com', 'www.nytimes.com', 'www.businessinsider.com', 'www.gfk.com', 'www.rugby.com', 'www.britannica.com', 'legallanguage.com', 'theledger.com', 'www.allmusic.com', 'iw.newsbank.com', 'www.nytimes.com', 'books.google.com', 'iw.newsbank.com', 'streetdirectory.com', 'www.mordorintelligence.com', 'www.statista.com', 'www.eulerhermes.com', 'www.foodnavigator.com', 'www.imdb.com', 'www.nature.com', 'in.reuters.com', 'www.britannica.com', 'query.nytimes.com', 'www.france-pub.com', 'books.google.com', 'www.time.com', 'books.google.com', 'www.fifa.com', 'www.smh.com', 'blog.hotelclub.com', 'edition.cnn.com', 'www.nationsencyclopedia.com', 'thetranslationcompany.com', 'www.theartnewspaper.com', 'www.britannica.com', 'www.statistiques-mondiales.com', 'www.franceway.com', 'www.la-croix.com', 'abcnews.go.com', 'www.ey.com', 'history.howstuffworks.com', 'observatoire.ojd.com', 'edition.cnn.com', 'www.bp.com', 'www.com', 'edition.cnn.com', 'www.businessweek.com', 'cannesguide.com', 'adherents.com', 'defense.com', 'books.google.com', 'www.paris-region.com', 'thetahititraveler.com', 'uk.franceguide.com', 'just-food.com', 'observatoire.ojd.com', 'books.google.com', 'books.google.com', 'www.lloydsbanktrade.com', 'nutraingredients.com', 'books.google.com', 'www.power-technology.com', 'books.google.com', 'www.statista.com', 'www.rfimusic.com', 'www.goodcooking.com', 'www.ifop.com', 'books.google.com', 'www.conventioncitoyenne.com', 'enotes.com', 'www.france24.com', 'topics.nytimes.com', 'www.etymonline.com', 'www.bbc.com', 'www.nytimes.com', 'www.fnsac-cgt.com', 'edition.cnn.com', 'books.google.com', 'www.smh.com', 'books.google.com', 'www.lecavalierbleu.com', 'www.france24.com', 'www.ojd.com', 'www.bbc.com', 'www.washingtonpost.com', 'www2.deloitte.com', 'iht.com', 'www.britannica.com', 'www.economist.com', 'www.bdpinternational.com', 'radiodramareviews.com', 'www.google.com', 'franceinlondon.com', 'climatechangepost.com', 'www.france24.com', 'books.google.com', 'dailyfinance.com', 'news.ambest.com', 'books.google.com', 'www.google.com', 'www.euractiv.com', 'www.uefa.com', 'www.nytimes.com', 'books.google.com', 'www.world-nuclear.org', 'www.coi-ioc.org', 'www.fao.org', 'www.eoearth.org', 'www.wto.org', 'www.lemans.org', 'www.ushmm.org', 'www.pewglobal.org', 'www.sipri.org', 'datatopics.worldbank.org', 'www.jstor.org', 'www.amnesty.org', 'ambafrance-us.org', 'www.ambafrance-dz.org', 'www.asylumineurope.org', 'whc.unesco.org', 'wayback.archive-it.org', 'www.un.org', 'transparency.org', 'www.ambafrance-ca.org', 'www.ctbto.org', 'understandfrance.org', 'unifrance.org', 'imf.org', 'www.un.org', 'loirevalley-worldheritage.org', 'stats.oecd.org', 'uis.unesco.org', 'www.indexoncensorship.org', 'www.ushmm.org', 'www.coi-ioc.org', 'www.pewglobal.org', 'data.oecd.org', 'www.unhcr.org', 'www.lemans.org', 'www.nobelprize.org', 'www.institutmontaigne.org', 'www.wto.org', 'humanistictexts.org', 'gesis.org', 'oecd-ilibrary.org', 'www.world-nuclear.org', 'www.pewglobal.org', 'hrw.org', 'www3.weforum.org', 'bigstory.ap.org', 'hosted.ap.org', 'data.worldbank.org', 'justfrance.org', 'wf-f.org', 'www.acs-aec.org', 'whc.unesco.org', 'www2.compareyourcountry.org', 'hdr.undp.org', 'www.globalreligiousfutures.org', 'obsarm.org', 'www.migrationpolicy.org', 'www.olympic.org', 'unstats.un.org', 'en.unesco.org', 'www.iea-pvps.org', 'unstats.un.org', 'www.migrationpolicy.org', 'www.world-nuclear.org', 'democracyweb.org', 'www.rpfrance-otan.org', 'www.ambafrance-cn.org', 'www.oecd.org', 'www.npr.org', 'www.wind-energy-the-facts.org', 'www.pewresearch.org', 'www.mathunion.org', 'www.indexoncensorship.org', 'www.weforum.org', 'oecdbetterlifeindex.org', 'ourworldindata.org', 'pris.iaea.org', 'www.hydropower.org', 'data.uis.unesco.org', 'hdr.undp.org', 'delegfrance-onu-geneve.org', 'www.npr.org', 'www.oecdbetterlifeindex.org', 'www.erudit.org', 'www.npr.org', 'ourworldindata.org', 'fas.org', 'www.iaea.org', 'www.oecd.org', 'www.francophonie.org', 'www.francophonie.org', 'www.nationalgallery.org', 'understandfrance.org', ['[[international affairs '], ['palgrave macmillan '], ['american journal of public health'], ['nature communications'], ['oxford university press'], ['transpl immunol. '], ['united nations world tourism organization ']]",5843419,Require autoconfirmed or confirmed access (no expiry set),350327,4 November 2001,63.224.38.xxx ,15836,33,2001-11-04,2001-11,2001
159,159,England,https://en.wikipedia.org/wiki/England,547,4,"['10.1098/rspb.2006.3627', '10.1080/02690940903166971', '10.1093/oxfordjournals.pubjof.a029948', '10.1038/1811754a0', '17002951', None, None, None, '1635457', None, None, None]","[['proceedings'], [' local economy'], ['publius'], ['nature ']]",42,64,0,82,0,14,342,0.07678244972577697,0.1170018281535649,0.14990859232175502,0.007312614259597806,0.0,0.20109689213893966,4,"['statistics.gov', 'www.gov', 'statistics.gov', 'www.gov', 'www.gov', 'ons.gov', 'www.ons.gov', 'statistics.gov', 'www.gov', 'www.ons.gov', 'ons.gov', 'www.culture.gov', 'number-10.gov', 'www.ons.gov', 'webarchive.nationalarchives.gov', 'www.ons.gov', 'www.ons.gov', 'royal.gov', 'www.gov', 'www.ons.gov', 'cabinetoffice.gov', 'webarchive.nationalarchives.gov', 'london.gov', 'www.gov', 'communities.gov', 'www.culture.gov', 'www.gov', 'www.gov', 'www.gov', 'www.dh.gov', 'www.gov', 'www.orr.gov', 'www.gov', 'www.ons.gov', 'cia.gov', 'www.gov', 'assets.publishing.service.gov', 'www.cia.gov', 'webarchive.nationalarchives.gov', 'nationalparks.gov', 'www.ons.gov', 'www.gov', 'royal.gov', 'statistics.gov', 'www.justice.gov', 'www.ons.gov', 'www.gov', 'statistics.gov', 'www.gov', 'www.hm-treasury.gov', 'cityoflondon.gov', 'webarchive.nationalarchives.gov', 'www.gov', 'www.metoffice.gov', 'www.gos.gov', 'www.dh.gov', 'webarchive.nationalarchives.gov', 'statistics.gov', 'homeoffice.gov', 'gos.gov', 'www.ons.gov', 'www.ons.gov', 'environment-agency.gov', 'www.gov', 'www.nytimes.com', 'online.wsj.com', 'sportbusiness.com', 'books.google.com', 'books.google.com', 'go.euromonitor.com', 'www.nytimes.com', 'www.theglobalist.com', 'books.google.com', 'www.newstatesman.com', 'galeon.com', 'books.google.com', 'www.worldatlas.com', 'statisticalyearbook11.ry.com', 'dictionary.law.com', 'money.uk.msn.com', 'www.renewableuk.com', 'www.renewableuk.com', 'www.ealingstudios.com', 'www.topuniversities.com', 'books.google.com', 'www.moorerail.com', 'www.britannica.com', 'www.medianewsline.com', 'economywatch.com', 'picturesofengland.com', 'www.powermag.com', 'books.google.com', 'spartacus-educational.com', 'www.cricinfo.com', 'www.fifa.com', 'www.users.waitrose.com', 'britainusa.com', 'fifa.com', 'facebook.com', 'www.medianewsline.com', 'travelsignposts.com', 'www.rolls-royce.com', 'eurotunnel.com', 'books.google.com', 'britannia.com', 'theculturetrip.com', 'visitbirmingham.com', 'dictionary.oed.com', 'books.google.com', 'britannica.com', 'rugbyfootballhistory.com', 'www.bloomberg.com', 'encarta.msn.com', 'edition.cnn.com', 'www.yaelf.com', 'findarticles.com', 'rankings.ft.com', 'history.com', 'bleacherreport.com', 'books.google.com', 'riaa.com', 'www.cricinfo.com', 'books.google.com', 'britannica.com', 'www.cincodias.com', 'books.google.com', 'books.google.com', 'www.time.com', 'www.pteducation.com', 'www.ppluk.com', 'metoffice.com', 'theworlds50best.com', 'books.google.com', 'heritage-key.com', 'dictionary.oed.com', 'www.americanheritage.com', 'worldsquash2008.com', 'britannica.com', 'artinfo.com', 'eitb24.com', 'www.newstatesman.com', 'books.google.com', 'www.etymonline.com', 'books.google.com', 'www.pgatour.com', 'www.dawn.com', 'www.bfi.org', 'www.english-heritage.org', 'www.churchofengland.org', 'www.royal-navy.org', 'www.summitpost.org', 'www.un.org', 'www.sciencemuseum.org', 'www.english-heritage.org', 'www.tate.org', 'www.geo-east.org', 'royalsociety.org', 'designatedsites.naturalengland.org', 'www.ihbc.org', 'www.thersa.org', 'www.instituteforgovernment.org', 'www.magakernow.org', 'www.goaldentimes.org', 'welshjournals.llgc.org', 'pdfs.semanticscholar.org', 'stone-circles.org', 'whc.unesco.org', 'www.nationaltrust.org', 'data.worldbank.org', 'britishmuseum.org', 'www.oecd.org', 'www.pbs.org', 'royalsociety.org', 'royalsociety.org', 'www.icons.org', 'pewresearch.org', 'www.rhs.org', 'designatedsites.naturalengland.org', 'www.iso.org', 'www.heroicage.org', 'www.cambridge.org', 'english-heritage.org', 'whc.unesco.org', 'royalsociety.org', 'www.artscouncil.org', 'www.nationaltrust.org', 'www.linguae-celticae.org', 'www.magakernow.org', ['proceedings'], [' local economy'], ['publius'], ['nature ']]",9316,Require administrator access (no expiry set),275583,17 October 2001,Zundark ,15044,6,2001-10-17,2001-10,2001
160,160,Gujarat,https://en.wikipedia.org/wiki/Gujarat,248,6,"['10.1890/i1540-9295-10-5-228', '10.1016/j.biocon.2011.02.009', '10.1080/00404969.2017.1294814', '10.1080/09614520050010214', '10.1023/b:bioc.0000040009.75090.8c', '10.1016/0024-6301(90)90104-c', None, None, None, None, None, None, None, None, None, None, None, None]","[['frontiers in ecology and the environment'], ['biological conservation '], ['textile history'], ['development in practice'], ['biodiversity '], ['long range planning ']]",19,18,0,147,0,0,58,0.07661290322580645,0.07258064516129033,0.592741935483871,0.024193548387096774,0.0,0.17338709677419356,6,"['soir.senate.ca.gov', 'www.nri.gujarat.gov', 'censusindia.gov', 'www.censusindia.gov', 'sycd.gov', 'agri.gujarat.gov', 'agri.gujarat.gov', 'censusindia.gov', 'gujsail.gujarat.gov', 'soir.senate.ca.gov', 'www.mospi.gov', 'gujsail.gujarat.gov', 'censusindia.gov', 'earthquake.usgs.gov', 'censusindia.gov', 'gujsail.gujarat.gov', 'planningcommission.gov', 'gujsail.gujarat.gov', 'tribune.com', 'www.dnaindia.com', 'books.google.com', 'books.google.com', 'www.nseindia.com', 'www.dnaindia.com', 'books.google.com', 'www.prosperity.com', 'books.google.com', 'books.google.com', 'books.google.com', 'articles.timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.hindustantimes.com', 'books.google.com', 'www.dnaindia.com', 'books.google.com', 'books.google.com', 'deshgujarat.com', 'www.financialexpress.com', 'tatasteel100.com', 'timesofindia.indiatimes.com', 'www.gujaratindia.com', 'gujaratindia.com', 'www.screenindia.com', 'books.google.com', 'www.thehindu.com', 'articles.timesofindia.indiatimes.com', 'rediff.com', 'books.google.com', 'www.moneycontrol.com', 'www.amul.com', 'economictimes.indiatimes.com', 'books.google.com', 'books.google.com', 'www.forbes.com', 'www.forbes.com', 'www.thehindubusinessline.com', 'culturopedia.com', 'books.google.com', 'books.google.com', 'www.firstpost.com', 'books.google.com', 'books.google.com', 'www.business-standard.com', 'mapsofindia.com', 'www.highbeam.com', 'articles.economictimes.indiatimes.com', 'books.google.com', 'www.indianexpress.com', 'cngcoins.com', 'www2.kenes.com', 'indianexpress.com', 'books.google.com', 'livemint.com', 'www.business-standard.com', 'indianexpress.com', 'indianexpress.com', 'theconversation.com', 'books.google.com', 'news.indiainfo.com', 'business-standard.com', 'books.google.com', 'www.forbes.com', 'books.google.com', 'gujaratirocks.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.gujaratindia.com', 'www.business-standard.com', 'books.google.com', 'newsonair.com', 'www.hindustantimes.com', 'www.britannica.com', 'books.google.com', 'gujaratindia.com', 'books.google.com', 'books.google.com', 'www.ndtv.com', 'deshgujarat.com', 'daily.bhaskar.com', 'books.google.com', 'www.bbc.com', 'economictimes.indiatimes.com', 'www.hindustantimes.com', 'books.google.com', 'www.amul.com', 'www.business-standard.com', 'books.google.com', 'www.time.com', 'the-south-asian.com', 'in.news.yahoo.com', 'books.google.com', 'www.ibnlive.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'deshgujarat.com', 'www.indianchristianity.com', 'articles.timesofindia.indiatimes.com', 'books.google.com', 'rbth.com', 'books.google.com', 'books.google.com', 'www.discoveredindia.com', 'timesofindia.indiatimes.com', 'www.gujaratindia.com', 'www.indianexpress.com', 'www.business-standard.com', 'books.google.com', 'www.hindustantimes.com', 'www.lonelyplanet.com', 'www.business-standard.com', 'articles.timesofindia.indiatimes.com', 'books.google.com', 'www.gujaratindia.com', 'rediff.com', 'books.google.com', 'books.google.com', 'articles.economictimes.indiatimes.com', 'books.google.com', 'livemint.com', 'www.thehindubusinessline.com', 'books.google.com', 'www.moneycontrol.com', 'www.india-seminar.com', 'mapsofindia.com', 'books.google.com', 'articles.timesofindia.indiatimes.com', 'books.google.com', 'wingsbirds.com', 'www.screenindia.com', 'indianexpress.com', 'www.japancentreatama.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'worldpopulationreview.com', 'books.google.com', 'in.news.yahoo.com', 'gujaratindia.com', 'www.in.kpmg.com', 'deshgujarat.com', 'timesofindia.indiatimes.com', 'rbth.com', 'www.fsi.org', 'iranicaonline.org', 'scity.org', 'aims.org', 'prsindia.org', 'www.downtoearth.org', 'www.ibiblio.org', 'globaldatalab.org', 'eadl.org', 'www.rbi.org', 'prsindia.org', 'hdi.globaldatalab.org', 'www.rajsaubhag.org', 'cadgog.org', 'cato.org', 'sindhology.org', 'www.gandhiashram.org', 'gksgujarat.org', 'www.gujaratcmfellowship.org', ['frontiers in ecology and the environment'], ['biological conservation '], ['textile history'], ['development in practice'], ['biodiversity '], ['long range planning ']]",53707,Require administrator access (no expiry set),201301,16 May 2002,PierreAbbat ,8762,34,2002-05-16,2002-05,2002
161,161,Chams,https://en.wikipedia.org/wiki/Chams,98,7,"['10.1080/14442210600965174', '10.4000/moussons.976', '10.1080/14672715.1988.10412580', '10.1371/journal.pone.0036437', '10.1038/ncomms5689', '10.1163/1878464x-01001001', '10.3406/arch.2013.4389', None, None, None, '22586471', '25137359', None, None, None, None, None, '3346718', '4143916', None, None]","[[' the asia pacific journal of anthropology ', ' the australian national university '], ['recherches en sciences sociales sur l', 'moussons '], [' ben kiernan', ' bulletin of concerned asian scholars '], ['plos one '], ['nature communications '], ['journal of islamic manuscripts'], ['archipel ']]",7,1,0,59,0,0,24,0.07142857142857142,0.01020408163265306,0.6020408163265306,0.07142857142857142,0.0,0.15306122448979592,7,"['state.gov', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'news.nationalgeographic.com', 'books.google.com', 'thailandsworld.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.nationalgeographic.com', 'books.google.com', 'books.google.com', 'www.aljazeera.com', 'books.google.com', 'books.google.com', 'chamunesco.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.aljazeera.com', 'www.chamtoday.com', 'mvslim.com', 'books.google.com', 'www.chamtoday.com', 'www.chamtoday.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.atimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'phnompenhpost.com', 'phnompenhpost.com', 'news.nationalgeographic.com', 'books.google.com', 'books.google.com', 'books.google.com', 'drive.google.com', 'books.google.com', 'chamtoday.com', 'books.google.com', 'books.google.com', 'themuslimvibe.com', 'books.google.com', 'books.google.com', 'everyculture.com', 'chamtoday.com', 'www.atlaswalisongo.com', 'www.laoamericansports.com', 'books.google.com', 'books.google.com', 'zh.wikisource.org', 'vietspring.org', 'worldmap.org', 'cambodianscholars.org', 'englishkyoto-seas.org', 'scriptsource.org', 'www.eurekalert.org', [' the asia pacific journal of anthropology ', ' the australian national university '], ['recherches en sciences sociales sur l', 'moussons '], [' ben kiernan', ' bulletin of concerned asian scholars '], ['plos one '], ['nature communications '], ['journal of islamic manuscripts'], ['archipel ']]",153025,Allow all users (no expiry set),75438,29 November 2002,65.184.35.217 ,1134,1,2002-11-29,2002-11,2002
162,162,West Bengal,https://en.wikipedia.org/wiki/West_Bengal,293,0,[],[],36,30,0,132,0,1,95,0.12286689419795221,0.10238907849829351,0.45051194539249145,0.0,0.0,0.22525597269624573,0,"['labourbureaunew.gov', 'tourism.gov', 'www.westbengaltourism.gov', 'censusindia.gov', 'censusindia.gov', 'www.censusindia.gov', 'darjeeling.gov', 'www.censusindia.gov', 'www.trai.gov', 'www.censusindia.gov', 'censusindia.gov', 'wb.gov', 'mhrd.gov', 'niti.gov', 'www.censusindia.gov', 'www.mospi.gov', 'kolkataporttrust.gov', 'niti.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'www.wbhealth.gov', 'censusindia.gov', 'www.westbengaltourism.gov', 'legislativebodiesinindia.gov', 'censusindia.gov', 'purulia.gov', 'www.censusindia.gov', 'www.naac.gov', 'niti.gov', 'www.censusindia.gov', 'www.telegraphindia.com', 'books.google.com', 'indianexpress.com', 'www.wbidc.com', 'books.google.com', 'www.contemporaryart-india.com', 'books.google.com', 'www.thehindu.com', 'www.financialexpress.com', 'books.google.com', 'www.moneycontrol.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thestatesman.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.business-standard.com', 'books.google.com', 'rediff.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.telegraphindia.com', 'amsglossary.allenpress.com', 'books.google.com', 'www.webindia123.com', 'books.google.com', 'timesfoundation.indiatimes.com', 'www.telegraphindia.com', 'books.google.com', 'www.thehindubusinessline.com', 'economictimes.indiatimes.com', 'swachhindia.ndtv.com', 'books.google.com', 'www.telegraphindia.com', 'm.economictimes.com', 'www.telegraphindia.com', 'www.thehindu.com', 'www.economist.com', 'books.google.com', 'timesofindia.indiatimes.com', 'economictimes.indiatimes.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'www.flonnet.com', 'www.voanews.com', 'economictimes.indiatimes.com', 'books.google.com', 'www.telegraphindia.com', 'www.thehindu.com', 'www.espncricinfo.com', 'books.google.com', 'www.thestatesman.com', 'longlivesoccer.com', 'timesofindia.indiatimes.com', 'books.google.com', 'bangalinet.com', 'books.google.com', 'rediff.com', 'www.financialexpress.com', 'www.bloombergquint.com', 'www.telegraphindia.com', 'www.newindianexpress.com', 'books.google.com', 'www.webel-india.com', 'www.outlookindia.com', 'www.financialexpress.com', 'books.google.com', 'www.thehansindia.com', 'books.google.com', 'www.telegraphindia.com', 'archive.indianexpress.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'www.telegraphindia.com', 'books.google.com', 'news.outlookindia.com', 'www.aljazeera.com', 'books.google.com', 'archives.cnn.com', 'books.google.com', 'books.google.com', 'books.google.com', 'centreforaviation.com', 'www.kolmetro.com', 'books.google.com', 'www.telegraphindia.com', 'www.thehindu.com', 'indianexpress.com', 'indianexpress.com', 'www.hindustantimes.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'economictimes.indiatimes.com', 'www.thehansindia.com', 'books.google.com', 'books.google.com', 'www.livemint.com', 'www.calcuttaweb.com', 'books.google.com', 'www.telegraphindia.com', 'books.google.com', 'www.educationobserver.com', 'books.google.com', 'books.google.com', 'timesofindia.com', 'indianexpress.com', 'thediplomat.com', 'books.google.com', 'www.telegraphindia.com', 'books.google.com', 'dw.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'fifa.com', 'www.business-standard.com', 'www.webindia123.com', 'rbidocs.rbi.org', 'en.banglapedia.org', 'www.ibef.org', 'rbi.org', 'hdr.undp.org', 'whc.unesco.org', 'en.banglapedia.org', 'www.fsi.org', 'www.nobelprize.org', 'www.undp.org', 'govdocs.aquake.org', 'en.banglapedia.org', 'irfca.org', 'whc.unesco.org', 'en.banglapedia.org', 'www.thewbuhs.org', 'www.futurehealthsystems.org', 'irfca.org', 'nobelprize.org', 'indiankanoon.org', 'www.ibef.org', 'en.banglapedia.org', 'lakdiva.org', 'www.satp.org', 'kolkata.china-consulate.org', 'library.la84.org', 'hdi.globaldatalab.org', 'en.banglapedia.org', 'whc.unesco.org', 'www.dospiwb.org', 'rchiips.org', 'www.downtoearth.org', 'www.rbi.org', 'en.banglapedia.org', 'rchiips.org', 'www.ibef.org']",34040,Require administrator access (no expiry set),199852,23 December 2001,Hagedis ,4461,27,2001-12-23,2001-12,2001
163,163,Mauritius,https://en.wikipedia.org/wiki/Mauritius,225,5,"['10.1126/science.295.5560.1683', '10.1353/jwh.2003.0026', '10.1038/s41467-020-19493-3', '10.1080/0023656x.2013.804268', '10.1215/9780822386919-011', '11872833', None, '33293507', None, None, None, None, '7723057', None, None]","[['science'], ['[[journal of world history'], ['nature communications'], ['labor history '], ['duke university press']]",81,6,0,52,0,4,78,0.36,0.02666666666666667,0.2311111111111111,0.022222222222222223,0.0,0.4088888888888889,5,"['www.sl.nsw.gov', 'www.cia.gov', '2009-2017.state.gov', 'biot.gov', 'www.cia.gov', 'www.nsb.gov', 'www.country-data.com', 'search.yahoo.com', 'www.passengerterminaltoday.com', '(www.dw.com', 'www.nytimes.com', 'www.mauritiusmag.com', 'books.google.com', 'www.thehindu.com', 'www.thehindu.com', 'www.geoffreyrobertson.com', 'knoema.com', 'www.lemauricien.com', 'www.reuters.com', 'www.bbc.com', 'www.nytimes.com', 'www.mauritiustimes.com', 'pcacases.com', 'www.lemauricien.com', 'mauritiusgovernment.com', 'www.movingthenationforward.com', 'www.mauritiustimes.com', 'www.economist.com', 'www.mauritiustimes.com', 'kreolmagazine.com', 'www.google.com', 'www.lemauricien.com', 'www.youtube.com', 'taxsummaries.pwc.com', 'www.forbes.com', 'www.intercontinentaltrust.com', 'country.eiu.com', 'thediplomat.com', 'www.lematinal.com', 'www.bbc.com', 'www.lemauricien.com', 'www.climatechangenews.com', 'www.afrol.com', 'www.france24.com', 'www.reuters.com', 'www.telegraphindia.com', 'pcacases.com', 'www.lematinal.com', 'www.internationalcuisine.com', 'news.yahoo.com', 'www.eiu.com', 'www.dtos-mu.com', 'www.roughguides.com', 'www.lemauricien.com', 'dw.com', 'www.bbc.com', 'www.realclearworld.com', 'books.google.com', 'statsmauritius.govmu.org', 'police.govmu.org', 'www.govmu.org', 'statsmauritius.govmu.org', 'files.pca-cpa.org', 'culture.govmu.org', 'www.edbmauritius.org', 'www.govmu.org', 'foreign.govmu.org', 'www.usip.org', 'www.un.org', 'pmo.govmu.org', 'www.fraserinstitute.org', 'www.refworld.org', 'culture.govmu.org', 'statsmauritius.govmu.org', 'foreign.govmu.org', 'www.project-syndicate.org', 'www.icj-cij.org', 'www.eisa.org', 'vintagemauritius.org', 'www.mauritian-wildlife.org', 'ministry-education.govmu.org', 'culture.govmu.org', 'www.imf.org', 'www.pewforum.org', 'www.wmf.org', 'hsumauritius.org', 'www.govmu.org', 'www.govmu.org', 'www.globalinnovationindex.org', 'files.pca-cpa.org', 'files.pca-cpa.org', 'whc.unesco.org', 'data.worldbank.org', 'www.mauritius.org', 'hsumauritius.org', 'www.heritage.org', 'www.govmu.org', 'culture.govmu.org', 'culture.govmu.org', 'statsmauritius.govmu.org', 'commons.wikimedia.org', 'mauritiusassembly.govmu.org', 'statsmauritius.govmu.org', 'www.govmu.org', 'www.eisa.org', 'www.eisa.org', 'www.edbmauritius.org', 'www.doingbusiness.org', 'mauritiusassembly.govmu.org', 'statsmauritius.govmu.org', 'www.mauritian-wildlife.org', 'foreign.govmu.org', 'hdr.undp.org', 'www.usip.org', 'www.govmu.org', 'president.govmu.org', 'www.eisa.org', 'mauritiusassembly.govmu.org', 'www.globalreligiousfutures.org', 'mauritiusassembly.govmu.org', 'www.fscmauritius.org', 'culture.govmu.org', 'www.earthtimes.org', 'president.govmu.org', 'npcs.govmu.org', 'datahelpdesk.worldbank.org', 'archive.chagossupport.org', 'www3.weforum.org', 'unctad.org', 'culture.govmu.org', 'www.govmu.org', 'pmo.govmu.org', 'visionofhumanity.org', 'www.icij.org', 'vintagemauritius.org', 'imf.org', 'statsmauritius.govmu.org', 'culture.govmu.org', 'tourism.govmu.org', ['science'], ['[[journal of world history'], ['nature communications'], ['labor history '], ['duke university press']]",19201,Require administrator access (no expiry set),158107,28 September 2001,Koyaanis Qatsi ,8888,17,2001-09-28,2001-09,2001
164,164,Morocco,https://en.wikipedia.org/wiki/Morocco,200,8,"['10.1038/s41467-020-19493-3', '10.1086/430073', '10.1038/35002501', '10.1007/s10531-015-1042-1', '10.1093/biosci/bix014', '10.1377/hlthaff.26.4.1009', '10.1080/13629390902747491', '33293507', '15791543', '10706275', None, '28608869', '17630444', None, '7723057', '1199377', None, None, '5451287', '2898512', None]","[['nature communications'], ['the american journal of human genetics '], ['nature'], ['biodiversity and conservation'], ['bioscience'], [' health affairs '], [' mediterranean politics ']]",42,13,0,75,0,0,62,0.21,0.065,0.375,0.04,0.0,0.315,7,"['www.defense.gov', 'cia.gov', 'www.cia.gov', '2009-2017.state.gov', 'www.pncl.gov', 'www.tourisme.gov', 'www.cia.gov', 'whitehouse.gov', '2009-2017.state.gov', 'www.cbs.gov', 'www.loc.gov', 'www.sgg.gov', 'export.gov', 'groups.yahoo.com', 'www.moroccoworldnews.com', 'books.google.com', 'www.worldtimeserver.com', 'www.nationsencyclopedia.com', 'www.statoids.com', 'www.nytimes.com', 'finance.yahoo.com', 'books.google.com', 'www.britannica.com', 'www.aljazeera.com', 'lavieeco.com', 'www.reuters.com', 'www.aljazeera.com', 'encarta.msn.com', 'www.britannica.com', 'pages.eiu.com', 'nuqudy.com', 'www.britannica.com', 'www.ethnologue.com', 'statoids.com', 'books.google.com', 'www.google.com', 'www.britannica.com', 'northafricapost.com', 'www.britannica.com', 'www.indexmundi.com', 'www.nytimes.com', 'support.microsoft.com', 'news.yahoo.com', 'assets.opencrs.com', 'books.google.com', 'www.google.com', 'www.afrol.com', 'www.aljazeera.com', 'www.wellesnet.com', 'www.bbc.com', 'www.reuters.com', 'www.aljazeera.com', 'www.nature.com', 'www.moroccoworldnews.com', 'morocco-berbertrips.com', 'www.latimes.com', 'about.com', 'books.google.com', 'fescooking.com', 'www.sudestada.com', 'soccernet.espn.go.com', 'encarta.msn.com', 'nuqudy.com', 'uk.encarta.msn.com', 'books.google.com', 'books.google.com', 'moroccobusinessnews.com', 'www.moroccoworldnews.com', 'www.newframe.com', 'www.britannica.com', 'bbc.com', 'www.aljazeera.com', 'news.vice.com', 'www.ictj.com', 'www.timesofisrael.com', 'books.google.com', 'books.google.com', 'www.google.com', 'www.nytimes.com', 'books.google.com', 'www.irishtimes.com', 'books.google.com', 'www.christianitytoday.com', 'knoema.com', 'books.google.com', 'maroccankitchenrecipes.blogspot.com', 'books.google.com', 'www.britannica.com', 'www.africanconservation.org', 'www.refworld.org', 'ccisabroad.org', 'minurso.unmissions.org', 'www.francophonie.org', 'read.oecd-ilibrary.org', 'www.bjpa.org', 'data.worldbank.org', 'www.amnestyusa.org', 'www.refworld.org', 'www.imf.org', 'memrieconomicblog.org', 'freedomhouse.org', 'hdr.undp.org', 'journals.plos.org', 'unesdoc.unesco.org', 'www.iso.org', 'www.icj.org', 'www.pewforum.org', 'data.worldbank.org', 'www.youthindex.org', 'migrationinformation.org', 'portal.unesco.org', 'data.worldbank.org', 'www.un.org', 'www.jewishvirtuallibrary.org', 'data.worldbank.org', 'www.francophonie.org', 'www.refworld.org', 'data.worldbank.org', 'data.worldbank.org', 'www.youthindex.org', 'www.hrw.org', 'www.realinstitutoelcano.org', 'www.afdb.org', 'jewishvirtuallibrary.org', 'www.migrationinformation.org', 'www.go-south.org', 'hrw.org', 'www.refworld.org', 'data.worldbank.org', 'www.un.org', ['nature communications'], ['the american journal of human genetics '], ['nature'], ['biodiversity and conservation'], ['bioscience'], [' health affairs '], [' mediterranean politics ']]",19291,Require administrator access (no expiry set),152966,23 May 2001,KoyaanisQatsi ,9141,9,2001-05-23,2001-05,2001
165,165,Genoa,https://en.wikipedia.org/wiki/Genoa,100,1,"['10.1093/acref/9780195130751.001.0001', None, None]",[['oxford university press ']],3,1,0,29,0,0,66,0.03,0.01,0.29,0.01,0.0,0.05,1,"['www.parliament.nsw.gov', 'portofinoworld.com', 'turismo.com', 'weather2travel.com', 'www.com', 'www.com', 'www.linkedin.com', 'books.google.com', 'books.google.com', 'www.embassypages.com', 'www.britannica.com', 'azerbaijans.com', 'ilsole24ore.com', 'www.crwflags.com', 'www.bloomberg.com', 'books.google.com', 'world66.com', 'www.nationsencyclopedia.com', 'www.britannica.com', 'www.com', 'moovitapp.com', 'books.google.com', 'books.google.com', 'www.com', 'moovitapp.com', 'www.linkedin.com', 'news.com', 'smart.com', 'www.ilsole24ore.com', 'www.britannica.com', 'data.un.org', 'www.connectedurbandevelopment.org', 'danielea.altervista.org', ['oxford university press ']]",47332321,Allow all users (no expiry set),124961,25 February 2002,151.24.145.xxx ,4046,3,2002-02-25,2002-02,2002
166,166,Tuscany,https://en.wikipedia.org/wiki/Tuscany,41,0,[],[],4,0,0,12,0,0,25,0.0975609756097561,0.0,0.2926829268292683,0.0,0.0,0.0975609756097561,0,"['books.google.com', 'books.google.com', 'books.google.com', 'about.com', 'books.google.com', 'books.google.com', 'go.euromonitor.com', 'books.google.com', 'books.google.com', 'travelguide.affordabletours.com', 'books.google.com', 'www.citemedmode.com', 'library.thinkquest.org', 'www.learner.org', 'hdi.globaldatalab.org', 'library.thinkquest.org']",21967242,Allow all users (no expiry set),57106,25 September 2001,213.140.9.xxx ,2384,11,2001-09-25,2001-09,2001
167,167,Portugal,https://en.wikipedia.org/wiki/Portugal,319,12,"['10.1038/s41467-020-19493-3', '10.1080/00437956.1979.11435671', '10.1017/s1574019606000812', '10.1007/s10531-004-5015-z', '10.1038/sdata.2016.91', '10.3406/rbph.1957.2022', '10.1007/s10531-016-1141-7', '10.1006/jmsc.2001.1060', '10.1111/j.1468-0289.2012.00658.x', '10.1093/biosci/bix014', '10.1086/513477', '10.14195/0872-0851_43_7', '33293507', None, None, None, '27727236', None, None, None, None, '28608869', '17436249', None, '7723057', None, None, None, '5058334', None, None, None, None, '5451287', '1852743', None]","[['nature communications'], ['word'], ['european constitutional law review'], ['biodiversity and conservation ', '[[springer science'], ['scientific data ', '[[nature '], ['revue belge de philologie et d'], ['biodiversity and conservation '], ['ices journal of marine science '], ['economic history review '], ['bioscience'], ['american journal of human genetics '], ['revista filosófica de coimbra ']]",32,8,0,85,0,1,181,0.10031347962382445,0.025078369905956112,0.2664576802507837,0.03761755485893417,0.0,0.16300940438871472,12,"['www.cia.gov', 'www.st.nmfs.noaa.gov', 'cia.gov', 'portugal.gov', 'www.mmc.gov', 'azores.gov', 'ibge.gov', 'cia.gov', 'books.google.com', 'algarvedailynews.com', 'www.reuters.com', 'www.theportugalnews.com', 'www.euromonitor.com', 'curiousread.com', 'www.euronews.com', 'eupedia.com', 'www.youtube.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.reuters.com', 'www.prison-insider.com', 'theportugalnews.com', 'liveandinvestoverseas.com', 'countryeconomy.com', 'mileniostadium.com', 'worldtravelawards.com', 'www.10best.com', 'globalgolfermag.com', 'www.nytimes.com', 'www.nytimes.com', 'www.devdiscourse.com', 'www.historyireland.com', 'history.com', 'www.totaltele.com', 'oilprice.com', 'books.google.com', 'khazaria.com', 'golisbon.com', 'okonomos.weebly.com', 'www.france24.com', 'books.google.com', 'eduardodias.com', 'countryeconomy.com', 'books.google.com', 'books.google.com', 'listafterlist.com', 'books.google.com', '2.deloitte.com', 'embaixada-portugal-brasil.blogspot.com', 'washingtonindependent.com', 'theportugalnews.com', 'www.time.com', 'www.topuniversities.com', 'economist.com', 'www.time.com', 'books.google.com', 'uk.reuters.com', 'books.google.com', 'www.eupedia.com', 'worldtravelawards.com', 'unrv.com', 'www.statista.com', 'www.britannica.com', 'uk.reuters.com', 'www.ekathimerini.com', 'whalewatchingazores.com', 'diarioeconomico.com', 'www.youtube.com', 'www.oed.com', 'economist.com', 'britannica.com', 'infoescola.com', 'www.travelpulse.com', 'www.europesun.com', 'notapositiva.com', 'tripwix.com', 'punchng.com', 'www.numbeo.com', 'etymonline.com', 'www.ft.com', 'www.statista.com', 'visitportugal.com', 'www.economist.com', 'tecmaia.com', 'worldtravelawards.com', 'www.ft.com', 'www.comunidadeculturaearte.com', 'theportugalnews.com', 'books.google.com', 'investingnews.com', 'books.google.com', 'www.scientificamerican.com', 'www.imf.org', 'prisonstudies.org', 'prisonstudies.org', 'data.worldbank.org', 'seatemperature.org', 'www.imf.org', 'www.oecd.org', 'stats.oecd.org', 'www.wdl.org', 'hdi.globaldatalab.org', 'globalbioclimatics.org', 'www.laphamsquarterly.org', 'www.worldcat.org', 'seatemperature.org', 'www.iea.org', 'data.oecd.org', 'jewishvirtuallibrary.org', 'ourworldindata.org', 'www.cato.org', 'imf.org', 'sinestecnopolo.org', 'hdr.undp.org', 'www.worldcat.org', 'worldcat.org', 'www.un.org', 'imf.org', 'ourworldindata.org', 'www.oecd.org', 'www.constituteproject.org', 'hdi.globaldatalab.org', 'www.fao.org', 'www.worldcat.org', ['nature communications'], ['word'], ['european constitutional law review'], ['biodiversity and conservation ', '[[springer science'], ['scientific data ', '[[nature '], ['revue belge de philologie et d'], ['biodiversity and conservation '], ['ices journal of marine science '], ['economic history review '], ['bioscience'], ['american journal of human genetics '], ['revista filosófica de coimbra ']]",23033,Require administrator access (no expiry set),291374,15 March 2001,Cdani ,20002,55,2001-03-15,2001-03,2001
168,168,Kathmandu,https://en.wikipedia.org/wiki/Kathmandu,131,4,"['10.3390/rs1030534', '10.1016/j.apgeog.2009.10.002', '10.1016/j.cities.2007.10.001', '10.1016/j.compenvurbsys.2010.07.005', None, None, None, None, None, None, None, None]","[['remote sensing'], ['applied geography'], ['cities'], ['computers']]",20,23,0,48,0,1,35,0.15267175572519084,0.17557251908396945,0.366412213740458,0.030534351145038167,0.0,0.35877862595419846,4,"['www.kathmandu.gov', 'www.kathmandu.gov', 'www.kathmandu.gov', 'www.kathmandu.gov', 'www.kathmandu.gov', 'kathmandu.gov', 'www.dhm.gov', 'pollution.gov', 'kathmandu.gov', 'www.kathmandu.gov', 'censusnepal.cbs.gov', 'www.kathmandu.gov', 'www.cia.gov', 'www.kathmandu.gov', 'www.kathmandu.gov', 'airnow.gov', 'www.kathmandu.gov', 'www.kathmandu.gov', 'www.kathmandu.gov', '2001-2009.state.gov', 'www.kathmandu.gov', 'cbs.gov', 'www.kathmandu.gov', 'asiatravel.com', 'books.google.com', 'chandragirihills.com', 'books.google.com', 'kathmandukingsxi.com', 'www.asiatravel.com', 'nepalitimes.com', 'thehimalayantimes.com', 'worldpopulationreview.com', 'www.nytimes.com', 'www.fifa.com', 'www.spacesnepal.com', 'routesonline.com', 'buddhim.20m.com', 'www.nepalitimes.com', 'www.nationalgeographic.com', 'katmandu-hotels.com', 'nepalnews.com', 'www.economist.com', 'nepalmandal.com', 'www.facebook.com', 'bossnepal.com', 'www.tripadvisor.com', 'nepalitimes.com', 'ekantipur.com', 'turkishairlines.com', 'archive.nepalitimes.com', 'ekantipur.com', 'docs.google.com', 'kathmandupost.com', 'thehimalayantimes.com', 'www.ekantipur.com', 'www.nepalitimes.com', 'www.nepalvista.com', 'thehimalayantimes.com', 'books.google.com', 'kathmandupost.com', 'www.healio.com', 'apostolicnunciatureindia.com', 'www.expeditionsnepal.com', 'visitnepal.com', 'www.newatravels.com', 'archive.nepalitimes.com', 'books.google.com', 'jwajalapa.com', 'kathmandupost.ekantipur.com', 'cpruscha.com', 'medchrome.com', 'www.caanepal.org', 'gorkhapatra.org', 'unesdoc.unesco.org', 'unesdoc.unesco.org', 'documents.worldbank.org', 'rmaf.org', 'unesco.org', 'nepalmap.org', 'www.fan.org', 'dsbcproject.org', 'www.princemahidolaward.org', 'jazzmandu.org', 'kathmanduarts.org', 'www.iied.org', 'www.globalbioclimatics.org', 'www.worldbank.org', 'www.therisingnepal.org', 'nepal.saarctourism.org', 'nepal.saarctourism.org', 'varghesepaul.org', ['remote sensing'], ['applied geography'], ['cities'], ['computers']]",17168,Allow all users (no expiry set),140219,6 November 2001,62.253.64.xxx ,4672,26,2001-11-06,2001-11,2001
169,169,Western culture,https://en.wikipedia.org/wiki/Western_culture,191,10,"['10.2307/2598327', '10.1017/s0022050700021100', '10.1038/053516a0', '10.2307/750865', '10.1191/0266355406gh380oa', '10.1111/1468-0289.00084', '10.1109/t-aiee.1942.5058456', '10.1080/14786441108564683', '10.2307/20029452', '10.2307/2707514', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None]","[['the economic history review '], ['journal of economic history '], ['nature '], ['journal of the warburg and courtauld institutes '], ['german history '], ['the economic history review '], ['transactions of the american institute of electrical engineers '], ['the london'], ['foreign affairs '], ['journal of the history of ideas ']]",18,7,0,34,0,1,121,0.09424083769633508,0.03664921465968586,0.17801047120418848,0.05235602094240838,0.0,0.18324607329842932,10,"['history.nasa.gov', 'state.gov', 'history.nasa.gov', 'www.jpl.nasa.gov', 'www.jpl.nasa.gov', 'www.nasa.gov', '2001-2009.state.gov', 'caselaw.lp.findlaw.com', 'books.google.com', 'actualitechretienne.files.wordpress.com', 'www.livinginternet.com', 'books.google.com', 'www.sciencedaily.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'books.google.com', 'www.timemaps.com', 'www.britannica.com', 'www.usatoday.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'britannica.com', 'www.nrbookservice.com', 'books.google.com', 'books.google.com', 'encarta.msn.com', 'www.britannica.com', 'www.oxforddictionaries.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'pewforum.org', 'www.worldcat.org', 'pewforum.org', 'minneapolisfed.org', 'pewforum.org', 'deirdremccloskey.org', 'broughttolife.sciencemuseum.org', 'www.sfmuseum.org', 'www.khanacademy.org', 'www.catholiceducation.org', 'minneapolisfed.org', 'pewforum.org', 'pewforum.org', 'www.bipm.org', 'www.fgi-tbff.org', 'usma.org', 'pewforum.org', 'plus.maths.org', ['the economic history review '], ['journal of economic history '], ['nature '], ['journal of the warburg and courtauld institutes '], ['german history '], ['the economic history review '], ['transactions of the american institute of electrical engineers '], ['the london'], ['foreign affairs '], ['journal of the history of ideas ']]",21208262,Allow all users (no expiry set),116793,18 January 2004,Gabbe ,4127,16,2004-01-18,2004-01,2004
170,170,China,https://en.wikipedia.org/wiki/China,697,25,"['10.1126/science.336.6080.402', '10.1017/jch.2017.45', '10.2307/2659525', '10.1017/s0003055413000014', '10.2307/2950087', '10.1787/9789264230040-en', '10.1111/j.1728-4457.2013.00555.x', '10.1086/681664', '10.1016/j.chieco.2018.10.010', '10.1177/186810261104000201', '10.1038/d41586-020-03402-1', '10.1073/pnas.1919850117', '10.1038/sdata.2018.214', '10.1080/10670564.2021.1893558', '10.22439/cjas.v35i1.5400', '10.3760/cma.j.issn.0254-6450.2020.02.003', '10.1126/science.acx9657', '10.1038/s41467-020-19493-3', '10.1093/heapro/dah105', '10.1162/016228805775124534', '10.1038/nature07741', '10.1016/j.quascirev.2013.06.030', '10.1007/s13524-017-0595-x', '10.1038/d41586-020-03165-9', '10.34667/tind.44315', '22539691', None, None, None, None, None, None, '31431804', None, None, '33262500', '32978301', '30375988', None, None, '32064853', '34793217', '33293507', '14976170', None, '19279636', None, '28762036', '33177687', None, None, None, None, None, None, None, None, '6701844', None, None, None, '7568317', '6207062', None, None, None, None, '7723057', None, None, None, None, None, None, None]","[[' science'], ['the journal of chinese history', '[[cambridge university press'], ['journal of asian studies'], ['american political science review'], ['[[the australian journal of chinese affairs'], ['[[organisation for economic co-operation and development'], ['[[population and development review'], ['[[the china journal'], ['[[china economic review '], ['journal of current chinese affairs'], ['nature'], ['[[proceedings of the national academy of sciences'], ['scientific data'], ['[[journal of contemporary china'], ['the copenhagen journal of asian studies', '[[copenhagen business school'], ['zhonghua liu xing bing xue za zhi ', 'zh'], ['science '], ['nature communications'], ['[[health promotion international'], ['[[international security '], ['nature'], ['[[quaternary science reviews'], ['[[demography '], ['nature'], ['world intellectual property organization']]",112,40,0,335,0,9,176,0.1606886657101865,0.05738880918220947,0.4806312769010043,0.035868005738880916,0.0,0.2539454806312769,25,"['en.cnta.gov', 'www.state.gov', 'www.eric.ed.gov', 'www.mas.gov', 'www.stats.gov', 'www.hkma.gov', 'www.cia.gov', 'www.cia.gov', 'www.stats.gov', 'loc.gov', 'en.moe.gov', 'environment.gov', 'www.defense.gov', 'www.nsf.gov', 'english.www.gov', 'lcweb2.loc.gov', 'ministers.treasury.gov', 'en.moe.gov', 'www.wenzhou.gov', 'www.nps.gov', 'www.sara.gov', 'en.moe.gov', 'www.cia.gov', 'www.cia.gov', 'www.nga.gov', 'moe.gov', 'www.nra.gov', 'en.moe.gov', 'www.usgs.gov', 'english.gov', 'nhfpc.gov', 'lcweb2.loc.gov', 'lcweb2.loc.gov', 'www.npc.gov', 'www.cia.gov', 'www.stats.gov', 'en.moe.gov', 'eric.ed.gov', 'www.gov', 'www.nsf.gov', 'mongabay.com', 'chinatoday.com', 'books.google.com', 'books.google.com', 'image101.360doc.com', 'www.nytimes.com', 'books.google.com', 'npcobserver.com', 'www.nytimes.com', 'books.google.com', 'www.nytimes.com', 'www.ft.com', 'articles.washingtonpost.com', 'smetimes.tradeindia.com', 'www.bbc.com', 'www.cnbc.com', 'www.bbc.com', 'books.google.com', 'www.nytimes.com', 'www.scmp.com', 'www.power-technology.com', 'www.chinafile.com', 'books.google.com', 'english.peopledaily.com', 'www.globalfirepower.com', 'www.nytimes.com', 'www.nytimes.com', 'www.taipeitimes.com', 'shanghairanking.com', 'news.xinhuanet.com', 'news.xinhuanet.com', 'www.spacedaily.com', 'nasaspaceflight.com', 'www.nytimes.com', 'www.csmonitor.com', 'books.google.com', 'www.power-technology.com', 'www.chinadaily.com', '360doc.com', 'time.com', 'www.nytimes.com', 'www.mobileworldlive.com', 'www.theodora.com', 'www.visualcapitalist.com', 'railway-technology.com', 'books.google.com', 'books.google.com', 'english.people.com', 'thestar.com', 'www.washingtonpost.com', 'www.britannica.com', 'www.washingtonpost.com', 'www.cnn.com', 'docin.com', 'cnnmoney.com', 'www.reuters.com', 'www.reuters.com', 'www.visualcapitalist.com', 'books.google.com', 'www.piie.com', 'www.forbes.com', 'dictionary.reference.com', 'www.nytimes.com', 'antpedia.com', 'www.reuters.com', 'books.google.com', 'apnews.myway.com', 'ceicdata.com', 'www.theodora.com', 'markets.businessinsider.com', 'www.wsj.com', 'img.webme.com', 'www.cnki.com', 'www.highbeam.com', 'books.google.com', 'www.ft.com', 'qz.com', 'd.wanfangdata.com', 'www.reuters.com', 'www.cnn.com', 'www.theglobeandmail.com', 'www.britannica.com', 'books.google.com', 'www.hollywoodreporter.com', 'www.nytimes.com', 'chinasportsbiz.com', 'www.bloomberg.com', 'www.mysinchew.com', 'www.economist.com', 'www.washingtonpost.com', 'www.aljazeera.com', 'www.mckinsey.com', 'www.theworldofchinese.com', 'www.aa.com', 'www.emarketer.com', 'www.economist.com', 'endata.com', 'www.nytimes.com', 'www.forbes.com', 'books.google.com', 'www.scmp.com', 'olympics.com', 'alphahistory.com', 'www.nytimes.com', 'www.bloomberg.com', 'technode.com', 'www.statista.com', 'www.skyscrapercenter.com', 'www.businessweek.com', 'img.webme.com', 'books.google.com', 'english.people.com', 'asia.nikkei.com', 'www.nytimes.com', 'www.scmp.com', 'www.time.com', 'books.google.com', 'www.ipsos.com', 'www.investopedia.com', 'www.ft.com', 'www.statista.com', 'jaynestars.com', 'www.nytimes.com', 'www.bbc.com', 'qz.com', 'www.dawn.com', 'www.theatlantic.com', 'books.google.com', 'www.wsj.com', 'www.reuters.com', 'books.google.com', 'wanfangdata.com', 'books.google.com', 'money.cnn.com', 'www.ft.com', 'www.afr.com', 'books.google.com', 'alphahistory.com', 'www.nbcnews.com', 'about.com', 'shanghairanking.com', 'mongabay.com', 'www.swift.com', 'www.bbc.com', 'www.cnbc.com', 'www.history.com', 'books.google.com', 'www.scmp.com', 'www.bloomberg.com', 'www.economist.com', 'www.economist.com', 'books.google.com', 'www.washingtonpost.com', 'www.nst.com', 'www.cnbc.com', 'www.pwccn.com', 'www.statista.com', 'www.ig.com', 'thediplomat.com', 'news.xinhuanet.com', 'books.google.com', 'www.ft.com', 'www.forbes.com', 'wenku.baidu.com', 'www.nytimes.com', 'www.nippon.com', 'www.ethnologue.com', 'www.reuters.com', 'www.bbc.com', 'www.scientificamerican.com', 'www.bloomberg.com', 'www.xinhuanet.com', 'www.business-standard.com', 'www.dw.com', 'chinatoday.com', 'www.reuters.com', 'www.technologyreview.com', 'www.economist.com', 'www.timeshighereducation.com', 'www.valuewalk.com', 'www.baotounews.com', 'seattletimes.com', 'english.people.com', 'global.chinadaily.com', 'books.google.com', 'www.zdnet.com', 'blogs.forbes.com', 'books.google.com', 'qz.com', 'world.time.com', 'www.theatlantic.com', 'www.britannica.com', 'www.usatoday.com', 'www.history.com', 'www.statista.com', 'deadline.com', 'www.nytimes.com', 'www.reuters.com', 'books.google.com', 'books.google.com', 'thediplomat.com', 'books.google.com', 'www.bbc.com', 'www.reuters.com', 'www.timeshighereducation.com', 'cultural-china.com', 'www.reuters.com', 'books.google.com', 'www.bloomberg.com', 'www.cnki.com', 'www.shanghairanking.com', 'cleantechnica.com', 'www.nytimes.com', 'www.bbc.com', 'www.dw.com', 'www.bloomberg.com', 'foreignpolicy.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'www.nytimes.com', 'news.google.com', 'www.cnn.com', 'www.scmp.com', 'demographia.com', 'www.forbes.com', 'www.oed.com', 'www.forbes.com', 'www.bloomberg.com', 'books.google.com', 'www.bbc.com', 'www.bbc.com', 'qz.com', 'books.google.com', 'www.ddtjournal.com', 'www.xinhuanet.com', 'www.atimes.com', 'books.google.com', 'ph.news.yahoo.com', 'www.forbes.com', 'www.businessweek.com', 'www.gbm.hsbc.com', 'www.ft.com', 'www.reuters.com', 'www.ft.com', 'books.google.com', 'qz.com', 'www.bbc.com', 'books.google.com', 'www.reuters.com', 'books.google.com', 'www.mobileworldlive.com', 'london2012.com', 'www.xinhuanet.com', 'www.nytimes.com', 'www.bloomberg.com', 'www.seattletimes.com', 'www.chinesecio.com', 'www.scmp.com', 'books.google.com', 'www.statista.com', 'www.britannica.com', 'www.cnn.com', 'www.csmonitor.com', 'asia.nikkei.com', 'www.visualcapitalist.com', 'www.thoughtco.com', 'www.wsj.com', 'www.oed.com', 'www.chinabankingnews.com', 'books.google.com', 'books.google.com', 'news.xinhuanet.com', 'www.wsj.com', 'e.hznews.com', 'www.cnn.com', 'www.britannica.com', 'www.statista.com', 'english.peopledaily.com', 'www.statista.com', '360doc.com', 'sports.sohu.com', 'www.forbes.com', 'www.washingtonpost.com', 'english.people.com', 'global.chinadaily.com', 'www.bloomberg.com', 'books.google.com', 'www.bbc.com', 'www.nytimes.com', 'www.statista.com', 'www.usnews.com', 'yicaiglobal.com', 'www.britannica.com', 'www.britannica.com', 'www.bbc.com', 'www.timeshighereducation.com', 'www.cbsnews.com', 'www.thenation.com', 'www.timeshighereducation.com', 'www.feer.com', 'www.ft.com', 'www.statista.com', 'mongabay.com', 'www.washingtonpost.com', 'books.google.com', 'www.bloomberg.com', 'theconversation.com', 'www.cnki.com', 'apnews.myway.com', 'factsanddetails.com', 'www.usatoday.com', 'www.forbes.com', 'books.google.com', 'www.nbcnews.com', 'books.google.com', 'fortune.com', 'www.bloomberg.com', 'eastday.com', '360doc.com', 'mongabay.com', 'www.slate.com', 'books.google.com', 'www.washingtonpost.com', 'blogs.forbes.com', 'www.nytimes.com', 'books.google.com', 'transcripts.cnn.com', 'www.forbes.com', 'www.nytimes.com', 'www.timeshighereducation.com', 'physicsworld.com', 'www.mnn.com', 'www.worldatlas.com', 'www.britannica.com', 'ideas.repec.org', 'www.iea.org', 'www.nobelprize.org', 'asme.org', 'www.policyreview.org', 'www.imf.org', 'www.prb.org', 'www.nobelprize.org', 'www.pewforum.org', 'www.fao.org', 'www.olympic.org', 'data.worldbank.org', 'cwur.org', 'chinapower.csis.org', 'www.refworld.org', 'www.oecd.org', 'www.wto.org', 'www.unmultimedia.org', 'www.weforum.org', 'hdr.undp.org', 'www.cfr.org', 'www.imf.org', 'www.un.org', 'www.china.org', 'www.awea.org', 'data.worldbank.org', 'data.worldbank.org', 'www.worldbank.org', 'www.irena.org', 'data.worldbank.org', 'www.worldshipping.org', 'www.sciencemag.org', 'www.instituteforenergyresearch.org', 'data.worldbank.org', 'www.weforum.org', 'unstats.un.org', 'cybergeo.revues.org', 'www.npr.org', 'globalreligiousfutures.org', 'data.worldbank.org', 'www.fao.org', 'www.imf.org', 'www.pewresearch.org', 'www.cfr.org', 'china.org', 'www.rsc.org', 'imf.org', 'stats.ioinformatics.org', 'www.chathamhouse.org', 'www.hrw.org', 'www.migrationpolicy.org', 'globaldiplomacyindex.lowyinstitute.org', 'whc.unesco.org', 'literature.org', 'chinapower.csis.org', 'www.wssinfo.org', 'www.asiabusinesscouncil.org', 'www.nobelprize.org', 'www.nber.org', 'datatopics.worldbank.org', 'www.efchina.org', 'data.worldbank.org', 'www.ucsusa.org', 'www.metmuseum.org', 'www.iucnredlist.org', 'www.unwto.org', 'www.constituteproject.org', 'icho-official.org', 'iza.org', 'www.worldbank.org', 'data.worldbank.org', 'www.china.org', 'www.unesco.org', 'www.china.org', 'www.un.org', 'www.monthlyreview.org', 'www.weforum.org', 'www.nbr.org', 'fas.org', 'www.ecosensorium.org', 'www.oecd.org', 'datatopics.worldbank.org', 'www.cis.org', 'www.iea-pvps.org', 'data.worldbank.org', 'nobelprize.org', 'www.iucnredlist.org', 'www.sipri.org', 'cybergeo.revues.org', 'www.pewforum.org', 'data.worldbank.org', 'data.worldbank.org', 'data.oecd.org', 'archive.archaeology.org', 'www.weforum.org', 'www.ilo.org', 'www.ibiblio.org', 'openknowledge.worldbank.org', 'www.globalslaveryindex.org', 'climateactiontracker.org', 'www.lowyinstitute.org', 'imo-official.org', 'data.worldbank.org', 'www.unicef.org', 'www.oecd.org', 'cato.org', 'www.sino-platonic.org', 'www.imf.org', 'www.mathunion.org', 'asean.org', 'nobelprize.org', 'ipho-unofficial.org', [' science'], ['the journal of chinese history', '[[cambridge university press'], ['journal of asian studies'], ['american political science review'], ['[[the australian journal of chinese affairs'], ['[[organisation for economic co-operation and development'], ['[[population and development review'], ['[[the china journal'], ['[[china economic review '], ['journal of current chinese affairs'], ['nature'], ['[[proceedings of the national academy of sciences'], ['scientific data'], ['[[journal of contemporary china'], ['the copenhagen journal of asian studies', '[[copenhagen business school'], ['zhonghua liu xing bing xue za zhi ', 'zh'], ['science '], ['nature communications'], ['[[health promotion international'], ['[[international security '], ['nature'], ['[[quaternary science reviews'], ['[[demography '], ['nature'], ['world intellectual property organization']]",5405,Require administrator access (no expiry set),348223,23 October 2001,63.192.137.xxx ,19194,57,2001-10-23,2001-10,2001
171,171,Finland,https://en.wikipedia.org/wiki/Finland,389,6,"['10.1093/biosci/bix014', '10.1787/20755120-table1', '10.1111/1467-9477.00048', '10.1016/s0140-6736(10)62187-3', '10.21542/gcsp.2018.13', '10.1038/s41467-020-19493-3', '28608869', None, None, '21496911', '30083543', '33293507', '5451287', None, None, None, '6062761', '7723057']","[['bioscience'], ['oecd ilibrary '], ['[[scandinavian political studies'], ['[[the lancet'], ['global cardiology science '], ['nature communications']]",42,7,0,66,0,2,266,0.10796915167095116,0.017994858611825194,0.16966580976863754,0.015424164524421594,0.0,0.14138817480719795,6,"['www.cia.gov', 'cia.gov', '2009-2017.state.gov', 'lcweb2.loc.gov', '2001-2009.state.gov', 'www.cia.gov', 'memory.loc.gov', 's3.amazonaws.com', 'www.lifeinlapland.com', 'new.visitfinland.com', 'time.com', 'www.economist.com', 'www.nytimes.com', 's3.amazonaws.com', 'www.wsj.com', 'www.nytimes.com', 'oasisoftheseas.com', 'books.google.com', 'finance.yahoo.com', 'trip101.com', 'books.google.com', 'expat-finland.com', 'royalcaribbeanpresscenter.com', 'artsandculture.google.com', 'www.jarvisydan.com', 'thelatinlibrary.com', 'www.mozartforum.com', 'medalspercapita.com', 'travelofinland.com', 'www.irishtimes.com', 'statista.com', 'thehockeynews.com', 'europe-cities.com', 'prosperity.com', 'tabblo.com', 'www.mozartforum.com', 'foreignpolicy.com', 'www.economist.com', 'www.nytimes.com', 'www.discoverthebaltic.com', 'newsfeed.time.com', 'musicfinland.com', 'theculturetrip.com', 'www.bbc.com', 'www.cnn.com', 'independenttravelcats.com', 'books.google.com', 'topuniversities.com', 'www.euronews.com', 'www.helsinki-airport.com', 'www.awardsandshows.com', 'archive.wikiwix.com', 'goldenglobes.com', 'www.geocities.com', 'memphismagazine.com', 'www.upi.com', 'www.wearethemighty.com', 'theculturetrip.com', 'www.nytimes.com', 'www.wsj.com', 'books.google.com', 'about.com', 'happiness-report.s3.amazonaws.com', 's3.amazonaws.com', 'fiba.com', 'books.google.com', 'www.focus-economics.com', 'theculturetrip.com', 'edition.cnn.com', 'books.google.com', 'www.ft.com', 'www.famouscampaigns.com', 'scholarshipsineurope.com', 'natowatch.org', 'www.councilwomenworldleaders.org', 'intelnews.org', 'www.weforum.org', 'www.imf.org', 'globalhealthfacts.org', 'norden.org', 'siteresources.worldbank.org', 'www.efnil.org', 'eurydice.org', 'newseum.org', 'www.unevoc.unesco.org', 'hdrstats.undp.org', 'stats.oecd.org', 'www.wan-ifra.org', 'www3.weforum.org', 'floorball.org', 'constituteproject.org', 'data.unicef.org', 'oecd.org', 'ich.unesco.org', 'www.un.org', 'www.amnesty.org', 'www3.weforum.org', 'hdr.undp.org', 'freedomhouse.org', 'natowatch.org', 'www.imf.org', 'www3.weforum.org', 'tuomioja.org', 'nobelprize.org', 'reports.weforum.org', 'pewforum.org', 'www.democracyranking.org', 'www.oecd.org', 'worldaudit.org', 'transparency.org', 'knowablemagazine.org', 'ourworldindata.org', 'doingbusiness.org', 'fundforpeace.org', 'www.heritage.org', ['bioscience'], ['oecd ilibrary '], ['[[scandinavian political studies'], ['[[the lancet'], ['global cardiology science '], ['nature communications']]",10577,Require administrator access (no expiry set),262124,8 September 2001,Koyaanis Qatsi ,14349,39,2001-09-08,2001-09,2001
172,172,Macedonia (Greece),https://en.wikipedia.org/wiki/Macedonia_(Greece),154,5,"['10.1086/ajs505193', '10.3167/001430003782266107', '10.1111/j.1467-8306.2007.00545.x', '10.4467/20834624sl.16.006.5152', '10.1017/s0079497x00013396', None, None, None, None, None, None, None, None, None, None]","[['[[american journal of archaeology'], ['european judaism'], ['annals of the association of american geographers '], ['studia linguistica universitatis iagellonicae cracoviensis '], ['proceedings of the prehistoric society ']]",12,2,0,37,0,0,98,0.07792207792207792,0.012987012987012988,0.24025974025974026,0.032467532467532464,0.0,0.12337662337662338,5,"['state.gov', '2009-2017.state.gov', 'www.myjewishlearning.com', 'www.fraport-greece.com', 'www.findarticles.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.ekathimerini.com', 'books.google.com', 'foreignpolicy.com', 'books.google.com', 'newrepublic.com', 'books.google.com', 'www.timesofisrael.com', 'books.google.com', 'www.lonelyplanet.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.etymonline.com', 'books.google.com', 'books.google.com', 'www.discovergreece.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.lonelyplanet.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'www.ekathimerini.com', 'www.freewebs.com', 'books.google.com', 'www.findarticles.com', 'www.balcanicaucaso.org', 'www.greekembassy.org', 'www.balcanicaucaso.org', 'www.promacedonia.org', 'whc.unesco.org', 'www.ushmm.org', 'www.doaks.org', 'www.promacedonia.org', 'www.osce.org', 'www.promacedonia.org', 'journals.openedition.org', 'journals.openedition.org', ['[[american journal of archaeology'], ['european judaism'], ['annals of the association of american geographers '], ['studia linguistica universitatis iagellonicae cracoviensis '], ['proceedings of the prehistoric society ']]",2741895,Allow all users (no expiry set),122794,8 May 2002,12.149.100.21 ,4519,1,2002-05-08,2002-05,2002
173,173,Kerala,https://en.wikipedia.org/wiki/Kerala,704,10,"['10.1016/0305-750x(96)00015-0', '10.11646/zootaxa.4985.3.5', '10.2307/2690896', '10.2307/2758883', '10.1017/s0007123412000178', '10.1093/heapol/15.1.103', '10.1007/bf02702224', '10.1086/356288', None, None, '34186802', None, None, None, '10731241', None, None, '19066487', None, None, None, None, None, None, None, None, None]","[['[[world development '], ['[[zootaxa'], ['mathematics magazine '], ['pacific affairs '], ['british journal of political science '], ['health policy and planning '], ['proc indian acad sci '], ['isis '], ['health physics ']]",51,50,0,439,0,0,154,0.07244318181818182,0.07102272727272728,0.6235795454545454,0.014204545454545454,0.0,0.15767045454545456,9,"['finance.kerala.gov', 'main.trai.gov', 'www.prd.kerala.gov', 'india.gov', 'rajbhavan.kerala.gov', 'kerala.gov', 'community.data.gov', 'sdgindiaindex.niti.gov', 'india.gov', 'www.archive.india.gov', 'ecostat.kerala.gov', 'main.trai.gov', 'www.kerala.gov', 'www.ecostat.kerala.gov', 'www.imd.gov', 'www.kerala.gov', 'www.censusindia.gov', 'www.forest.kerala.gov', 'dhs.kerala.gov', 'kerala.gov', 'keralacm.gov', 'www.keralapwd.gov', 'kite.kerala.gov', 'www.censusindia.gov', 'india.gov', 'www.kerala.gov', 'ildm.kerala.gov', 'www.keralapwd.gov', 'www.keralapwd.gov', 'planningcommission.gov', 'censusindia.gov', 'spb.kerala.gov', 'dmg.kerala.gov', 'www.ecostat.kerala.gov', 'kerala.gov', 'mohua.gov', 'spb.kerala.gov', 'www.censusindia.gov', 'planningcommission.gov', 'www.prd.kerala.gov', 'mahe.gov', 'www.censusindia.gov', 'www.ecostat.kerala.gov', 'www.mospi.gov', 'www.censusindia.gov', 'archive.india.gov', 'legislative.gov', 'fisheries.kerala.gov', 'sametham.kite.kerala.gov', 'www.keralapwd.gov', 'www.thehindubusinessline.com', 'books.google.com', 'm.timesofindia.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'economictimes.indiatimes.com', 'thehindu.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'news.google.com', 'www.indianexpress.com', 'www.ndtv.com', 'www.newindianexpress.com', 'books.google.com', 'www.dnaindia.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'yentha.com', 'www.thehindu.com', 'www.thehindu.com', 'www.indushealthplus.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.mathrubhumi.com', 'www.tripays.com', 'www.indianexpress.com', 'www.indianmirror.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'm.timesofindia.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.business-standard.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'upscguide.com', 'www.thenewsminute.com', 'books.google.com', 'books.google.com', 'books.google.com', 'forbesindia.com', 'www.thehindu.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'timesofindia.indiatimes.com', 'economictimes.indiatimes.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.cnn.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'sports.ndtv.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'books.google.com', 'khelnow.com', 'www.the-aiff.com', 'www.financialexpress.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'www.thehindu.com', 'www.thehindu.com', 'books.google.com', 'english.manoramaonline.com', 'articles.timesofindia.indiatimes.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'www.rediff.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'rediff.com', 'www.thehindu.com', 'indianexpress.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'keralartc.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'www.thehindu.com', 'www.thehindu.com', 'books.google.com', 'www.arabnews.com', 'books.google.com', 'english.mathrubhumi.com', 'books.google.com', 'ibnlive.in.com', 'www.hindu.com', 'books.google.com', 'www.firstpost.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'keralaliterature.com', 'timesofindia.indiatimes.com', 'www.keralartc.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'in.finance.yahoo.com', 'books.google.com', 'google.com', 'timesofindia.indiatimes.com', 'www.hindu.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'articles.timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'www.khaleejtimes.com', 'www.thehindu.com', 'books.google.com', 'www.hindu.com', 'zeenews.india.com', 'books.google.com', 'www.thehindubusinessline.com', 'books.google.com', 'books.google.com', 'query.nytimes.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'biblestudytools.com', 'books.google.com', 'books.google.com', 'www.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'economictimes.indiatimes.com', 'www.onmanorama.com', 'www.mathrubhumi.com', 'books.google.com', 'www.hindu.com', 'books.google.com', 'www.hindu.com', 'indianexpress.com', 'articles.economictimes.indiatimes.com', 'www.thehindu.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'pravasikairali.com', 'www.livemint.com', 'www.hindu.com', 'www.bbc.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.ndtv.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'www.ndtv.com', 'www.hindu.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'dictionary.reference.com', 'books.google.com', 'www.hindu.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.onmanorama.com', 'www.hindu.com', 'books.google.com', 'books.google.com', 'dhsprogram.com', 'books.google.com', 'www.thehindu.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'www.asianage.com', 'economictimes.indiatimes.com', 'books.google.com', 'www.financialexpress.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.thehindubusinessline.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.hindu.com', 'books.google.com', 'www.outlookindia.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.youtube.com', 'books.google.com', 'books.google.com', 'the-aiff.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.rediff.com', 'economictimes.indiatimes.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'monstersandcritics.com', 'books.google.com', 'www.youtube.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'www.newindianexpress.com', 'www.thehindu.com', 'www.thehindu.com', 'www.business-standard.com', 'www.thehindu.com', 'books.google.com', 'www.madhyamam.com', 'books.google.com', 'www.dnaindia.com', 'books.google.com', 'www.thehindubusinessline.com', 'books.google.com', 'books.google.com', 'khsrcl.com', 'www.hindu.com', 'books.google.com', 'books.google.com', 'www.firstpost.com', 'books.google.com', 'books.google.com', 'www.deccanherald.com', 'www.mathrubhumi.com', 'www.thehindu.com', 'bbc.com', 'books.google.com', 'books.google.com', 'books.google.com', 'google.com', 'www.hindu.com', 'books.google.com', 'www.thehindu.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'nilamburnews.com', 'onlinestore.dcbooks.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.thehindu.com', 'www.hindu.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.newindianexpress.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'malayalam.news18.com', 'books.google.com', 'books.google.com', 'www.jagranjosh.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'english.mathrubhumi.com', 'books.google.com', 'www.thehindubusinessline.com', 'www.indianexpress.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.google.com', 'www.thehindu.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'slbckerala.com', 'afaqs.com', 'www.hindu.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'www.deccanchronicle.com', 'books.google.com', 'books.google.com', 'www.alstom.com', 'books.google.com', 'books.google.com', 'sportstar.thehindu.com', 'books.google.com', 'books.google.com', 'www.thehindubusinessline.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.hindu.com', 'books.google.com', 'www.newindianexpress.com', 'www.moneycontrol.com', 'books.google.com', 'www.travelportalofindia.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'www.rbi.org', 'threatenedtaxa.org', 'rchiips.org', 'www.cartage.org', 'ideas.repec.org', 'www.in.undp.org', 'rainforestinfo.org', 'www.ibef.org', 'www.corporationoftrivandrum.org', 'niyamasabha.org', 'www.keralatourism.org', 'niyamasabha.org', 'www.keralatourism.org', 'www.ncscm.org', 'www.kilaonline.org', 'www.keralatourism.org', 'www.gutenberg.org', 'keralaathletics.org', 'krpcds.org', 'rchiips.org', 'www.unesco.org', 'www.keralatourism.org', 'www.im4change.org', 'www.keralatourism.org', 'transparencyindia.org', 'www.kilaonline.org', 'www.ksudp.org', 'archive.transparency.org', 'krpcds.org', 'rbidocs.rbi.org', 'www.keralait.org', 'hdr.undp.org', 'www.unwire.org', 'www.keralatourism.org', 'www.ceped.org', 'churchmissionsociety.org', 'keralatourism.org', 'www.allindiajudges.org', 'www.keralatourism.org', 'churchmissionsociety.org', 'services.iriskf.org', 'www.keralatourism.org', 'siamese-heritage.org', 'hdi.globaldatalab.org', 'www.sruti.org', 'hdr.undp.org', 'www.ksidc.org', 'www.keralatourism.org', 'www.ncscm.org', 'www.trainweb.org', 'www.corporationoftrivandrum.org', ['[[world development '], ['[[zootaxa'], ['mathematics magazine '], ['pacific affairs '], ['british journal of political science '], ['health policy and planning '], ['proc indian acad sci '], ['isis '], ['health physics ']]",4349459,Require autoconfirmed or confirmed access (no expiry set),362953,31 October 2001,Ramesh ,15963,11,2001-10-31,2001-10,2001
174,174,Mongolia,https://en.wikipedia.org/wiki/Mongolia,145,4,"['10.1080/17441730902992067', '10.1038/s41467-020-19493-3', '10.3390/economies7020051', '10.1057/palgrave.fp.8200087', None, '33293507', None, None, None, '7723057', None, None]","[['asian population studies '], ['nature communications'], ['economies '], ['french politics ']]",26,10,0,40,0,1,64,0.1793103448275862,0.06896551724137931,0.27586206896551724,0.027586206896551724,0.0,0.27586206896551724,4,"['state.gov', 'www.cia.gov', 'gec.gov', '2009-2017.state.gov', 'www.cia.gov', 'mongolia.usembassy.gov', 'www.census.gov', 'www.loc.gov', 'www.loc.gov', 'dfat.gov', 'www.reuters.com', 'edition.cnn.com', 'www.upi.com', 'www.lodimapress.com', 'www.iht.com', 'www.britannica.com', 'www.britannica.com', 'www.ft.com', 'www.washingtonpost.com', 'www.britannica.com', 'asianart.com', 'www.scribd.com', 'infomongolia.com', 'mad-mongolia.com', 'www.pressreference.com', 'www.chriskaplonski.com', 'temperature.com', 'lonelyplanet.com', 'books.google.com', 'www.smh.com', 'www.economist.com', 'www.orientmag.com', 'books.google.com', 'www.businessinsider.com', 'books.google.com', 'www.economist.com', 'encyclopedia2.thefreedictionary.com', 'www.efinancialnews.com', 'news.nationalgeographic.com', 'www.pressreader.com', 'books.google.com', 'embassypages.com', 'www.e-mongol.com', 'www.bbc.com', 'mongolia-attractions.com', 'www.wunderground.com', 'books.google.com', 'thediplomat.com', 'thediplomat.com', 'www.worldpoliticsreview.com', 'www.jamestown.org', 'www.ocasia.org', 'rsf.org', 'churchofjesuschrist.org', 'blogs.adb.org', 'developmentprogress.org', 'www.unescap.org', 'www.wilsoncenter.org', 'freedomhouse.org', 'hdr.undp.org', 'www.jamestown.org', 'en.rsf.org', 'workspace.unpan.org', 'adventistyearbook.org', 'imf.org', 'www.bitig.org', 'www.fao.org', 'un.org', 'www.globalpolicy.org', 'hdr.undp.org', 'www.constitutionnet.org', 'data.worldbank.org', 'www.un.org', 'data.worldbank.org', 'www.issf-shooting.org', 'www.un.org', ['asian population studies '], ['nature communications'], ['economies '], ['french politics ']]",19271,Require administrator access (no expiry set),134321,23 May 2001,KoyaanisQatsi ,5969,1,2001-05-23,2001-05,2001
175,175,Fast food,https://en.wikipedia.org/wiki/Fast_food,92,20,"['10.1146/annurev.publhealth.22.1.309', '10.2105/ajph.2013.301677', '10.1001/jamapediatrics.2014.140', '10.1007/s00125-014-3382-x', '10.1111/nure.12031', '10.1371/journal.pone.0103543', '10.1525/gfc.2001.1.1.36', '10.1177/0009922814561742', '10.1111/j.1467-8594.2008.00322.x', '10.2307/3097205', '10.1016/j.nutres.2010.07.002', '10.1186/1479-5868-3-2', '10.1016/j.orcp.2008.03.004', '10.1155/2012/597924', '10.1016/j.appet.2016.11.016', '10.1093/ajcn/85.1.201', '10.1111/j.1748-720x.2007.00120.x', '10.1161/circulationaha.112.115923', '10.1108/01425450610683627', '10.1111/obr.12107', '11274524', '24625145', '24686476', '25303998', '23590707', '25062277', None, '25480321', None, None, '20851306', '16436207', '24351729', '22619703', '27864073', '17209197', '17341224', '22753305', None, '24102801', None, '3987573', None, '4221538', None, '4111613', None, None, None, None, None, '1397859', None, '3352603', None, None, None, '3401093', None, None]","[['annual review of public health'], [' american journal of public health'], ['[[jama pediatrics'], ['diabetologia'], ['nutrition reviews '], ['plos one'], ['gastronomica'], [' clinical pediatrics '], ['business and society review'], ['social problems'], ['nutrition research'], ['international journal of behavioral nutrition and physical activity'], ['obesity research '], [' journal of obesity '], ['appetite'], ['the american journal of clinical nutrition'], [' journal of law'], ['circulation'], ['employee relations'], ['obesity reviews ']]",12,2,0,25,0,2,31,0.13043478260869565,0.021739130434782608,0.2717391304347826,0.21739130434782608,0.0,0.3695652173913043,20,"['files.eric.ed.gov', 'bls.gov', 'www.franchisehelp.com', 'www.wienerwald.com', 'jpfarrell.blogspot.com', 'books.google.com', 'www.subway.com', 'www.globenewswire.com', 'www.burgerking.com', 'www.kfc.com', 'www.businessinsider.com', 'articles.latimes.com', 'www.livestrong.com', 'well.blogs.nytimes.com', 'parenting.blogs.nytimes.com', 'www.upi.com', 'www.eapplicants.com', 'www.vacationsmadeeasy.com', 'www.reuters.com', 'www.subway.com', 'www.nytimes.com', 'blogs.reuters.com', 'www.healthline.com', 'www.yum.com', 'www.wienerwald.com', 'franchisehelp.com', 'www.tacobell.com', 'pediatrics.aappublications.org', 'nelp.org', 'coloncancerfoundation.org', 'www.restaurant.org', 'uconnruddcenter.org', 'www.eurekalert.org', 'www.npr.org', 'www.yaleruddcenter.org', 'www.fastfoodmarketing.org', 'content.healthaffairs.org', 'www.cabdirect.org', 'ourlife.org', ['annual review of public health'], [' american journal of public health'], ['[[jama pediatrics'], ['diabetologia'], ['nutrition reviews '], ['plos one'], ['gastronomica'], [' clinical pediatrics '], ['business and society review'], ['social problems'], ['nutrition research'], ['international journal of behavioral nutrition and physical activity'], ['obesity research '], [' journal of obesity '], ['appetite'], ['the american journal of clinical nutrition'], [' journal of law'], ['circulation'], ['employee relations'], ['obesity reviews ']]",360101,Require autoconfirmed or confirmed access (no expiry set),58028,28 March 2002,Ed Poor ,5302,0,2002-03-28,2002-03,2002
176,176,Slovakia,https://en.wikipedia.org/wiki/Slovakia,162,4,"['10.1038/s41467-020-19493-3', '10.1080/09654310600852639', '10.1080/00438243.1978.9979728', '10.1093/biosci/bix014', '33293507', None, None, '28608869', '7723057', None, None, '5451287']","[['nature communications'], ['european planning studies '], ['world archaeology'], ['bioscience']]",20,8,0,27,0,2,102,0.12345679012345678,0.04938271604938271,0.16666666666666666,0.024691358024691357,0.0,0.19753086419753085,4,"['upn.gov', 'www.cia.gov', 'state.gov', 'lcweb2.loc.gov', 'www.cia.gov', '2009-2017.state.gov', 'www.loc.gov', 'www.cia.gov', 'slovakiasite.com', 'www.pressreleasepoint.com', 'www.aljazeera.com', 'books.google.com', 'slovakiasite.com', 'iihf.com', 'www.eset.com', 'www.ceeol.com', 'dictionary.reference.com', 'books.google.com', 'www.gallup.com', 'www.economist.com', 'books.google.com', 'iihf.com', 'industryweek.com', 'concise.britannica.com', 'wordpress.com', 'slovakiasite.com', 'books.google.com', 'www.slovensko.com', 'books.google.com', 'www.bloomberg.com', 'ta3.com', 'theconversation.com', 'books.google.com', 'mertsahinoglu.com', 'www.henleyglobal.com', 'www.oecd.org', 'slovakia.org', 'www.cybertruffle.org', 'www.worldcat.org', 'www.un.org', 'un.org', 'www.worldcat.org', 'www.slovakia.org', 'communistcrimes.org', 'wayback.archive-it.org', 'whc.unesco.org', 'hdr.undp.org', 'www.worldcat.org', 'communistcrimes.org', 'www.euforbih.org', 'imf.org', 'www.slovak-jewish-heritage.org', 'www.oecd.org', 'stats.oecd.org', 'web.worldbank.org', ['nature communications'], ['european planning studies '], ['world archaeology'], ['bioscience']]",26830,Require administrator access (no expiry set),153448,24 March 2001,Rob Salzman ,7796,9,2001-03-24,2001-03,2001
177,177,Amhara people,https://en.wikipedia.org/wiki/Amhara_people,139,12,"['10.1353/nas.2005.0004', 'abs/10.1080/14725840802417943', '10.1111/j.1749-6632.1962.tb50145.x', '10.1093/mq/lxi.1.47', '10.1017/hia.2016.13', '10.1093/afraf/adaa029', '10.2307/1158345', '10.1080/14725840802417943', '10.3406/ethio.2013.1539', '10.1111/j.1755-618x.1974.tb00004.x', '10.1163/18177565-90000138', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None]","[['northeast african studies'], ['african identities '], ['annals of the new york academy of sciences ', 'wiley-blackwell '], [' the musical quarterly '], ['history in africa'], ['african affairs'], ['africa ', 'cambridge university press  '], ['african identities'], ['annales d'], ['canadian review of sociology ', 'wiley-blackwell '], ['scrinium']]",10,2,0,46,0,1,68,0.07194244604316546,0.014388489208633094,0.33093525179856115,0.08633093525179857,0.0,0.17266187050359713,11,"['www.csa.gov', 'www.border.gov', 'books.google.com', 'books.google.com', 'www.google.com', 'www.ethnologue.com', 'addisstandard.com', 'www.ethiomedia.com', 'explorepartsunknown.com', 'books.google.com', 'www.britannica.com', 'www.brilliant-ethiopia.com', 'books.google.com', 'books.google.com', 'www.ethiopianreview.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'www.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.amharictube.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.ethiopianstories.com', 'books.google.com', 'writteninmusic.com', 'www.google.com', 'books.google.com', 'www.ethnologue.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.ethiopia-insight.com', 'www.ethnologue.com', 'books.google.com', 'books.google.com', 'www.africanews.com', 'www.britannica.com', 'ethiopiaforums.com', 'books.google.com', 'www.worldcat.org', 'npr.org', 'www.worldcat.org', 'www.worldcat.org', 'www.jstor.org', 'www.afropop.org', 'www.worldcat.org', 'catalog.ihsn.org', 'www.worldcat.org', 'www.senamirmir.org', ['northeast african studies'], ['african identities '], ['annals of the new york academy of sciences ', 'wiley-blackwell '], [' the musical quarterly '], ['history in africa'], ['african affairs'], ['africa ', 'cambridge university press  '], ['african identities'], ['annales d'], ['canadian review of sociology ', 'wiley-blackwell '], ['scrinium']]",355173,Allow all users (no expiry set),72570,2 November 2003,Bogdangiusca ,3196,38,2003-11-02,2003-11,2003
178,178,Byzantine Empire,https://en.wikipedia.org/wiki/Byzantine_Empire,484,29,"['10.2307/310399', '10.1017/s0034412500009094', '10.1093/past/84.1.3', '10.2307/2853672', '10.2307/1291170', '10.1093/ehr/xxvii.cvi.287', '10.3390/land7040153', '10.1080/00033798500200131', '10.12681/byzsym.857', '10.2307/1291127', '10.12681/byzsym.649', '10.2307/3168653', '10.2307/626864', '10.2307/294410', '10.2307/3591389', '10.7767/zrgka.1943.32.1.509', '10.2307/500639', '10.1017/s0362152900008722', '10.1007/bf02898434', '10.2307/624442', '10.1017/s0022050700096947', '10.1163/1568520991201687', '10.1177/03058298060340030201', '10.2307/1291256', '10.1086/486406', '10.1086/355661', '10.3828/978-0-85323-106-6', '10.1093/ehr/xc.ccclvii.721', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None]","[['harvard studies in classical philology '], ['religious studies '], ['past and present '], ['speculum '], ['dumbarton oaks papers '], ['the english historical review '], ['land ', 'mdpi ag '], ['annals of science '], ['byzantina symmeikta '], ['dumbarton oaks papers '], ['byzantina symmeikta '], ['church history '], ['the journal of hellenic studies '], ['the american journal of philology '], ['dumbarton oaks papers '], ['zeitschrift der savigny-stiftung für rechtsgeschichte'], ['american journal of archaeology '], ['tradition '], ['international journal of the classical tradition '], ['the journal of hellenic studies '], ['the journal of economic history '], ['journal of the economic and social history of the orient '], ['millennium'], ['dumbarton oaks papers '], ['the journal of religion '], ['[[isis ', (' astronomical works of gregory chioniades', ' chioniades', 'chioniades', 'v')], ['liverpool university press '], ['the english historical review ']]",17,0,0,40,0,0,398,0.03512396694214876,0.0,0.08264462809917356,0.05991735537190083,0.0,0.09504132231404959,28,"['books.google.com', 'www.lowtechmagazine.com', 'articles.latimes.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'concise.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.intratext.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.intratext.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'rbedrosian.com', 'denysmontandon.com', 'www.britannica.com', 'www.historytoday.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'www.doaks.org', 'www.doaks.org', 'www.worldhistory.org', 'www.worldhistory.org', 'www.ccel.org', 'www.metmuseum.org', 'www.doaks.org', 'www.romanity.org', 'www.worldcat.org', 'www.doaks.org', 'www.doaks.org', 'www.doaks.org', 'www.ams.org', 'www.worldcat.org', 'www.worldhistory.org', 'www.newadvent.org', 'www.jstor.org', ['harvard studies in classical philology '], ['religious studies '], ['past and present '], ['speculum '], ['dumbarton oaks papers '], ['the english historical review '], ['land ', 'mdpi ag '], ['annals of science '], ['byzantina symmeikta '], ['dumbarton oaks papers '], ['byzantina symmeikta '], ['church history '], ['the journal of hellenic studies '], ['the american journal of philology '], ['dumbarton oaks papers '], ['zeitschrift der savigny-stiftung für rechtsgeschichte'], ['american journal of archaeology '], ['tradition '], ['international journal of the classical tradition '], ['the journal of hellenic studies '], ['the journal of economic history '], ['journal of the economic and social history of the orient '], ['millennium'], ['dumbarton oaks papers '], ['the journal of religion '], ['[[isis ', (' astronomical works of gregory chioniades', ' chioniades', 'chioniades', 'v')], ['liverpool university press '], ['the english historical review ']]",16972981,Allow all users (no expiry set),233368,4 October 2001,MichaelTinkler ,12429,41,2001-10-04,2001-10,2001
179,179,Croatia,https://en.wikipedia.org/wiki/Croatia,317,8,"['10.1093/biosci/bix014', '10.18111/wtobarometereng.2019.17.1.2', '10.1093/oxfordjournals.ejil.a035834', '10.3935/rsp.v10i2.124', '10.1080/1462352032000149495', None, '10.1038/s41467-020-19493-3', '10.15291/geoadria.45', '28608869', None, None, None, None, '21682056', '33293507', None, '5451287', None, None, None, None, None, '7723057', None]","[['bioscience'], ['unwto world tourism barometer '], ['european journal of international law'], ['revija za socijalnu politiku'], ['[[journal of genocide research'], ['acta medico-historica adriatica', 'hrvatsko znanstveno društvo za povijest zdravstvene kulture'], ['nature communications'], ['geoadria', 'hrvatsko geografsko društvo ']]",23,10,0,69,0,0,208,0.07255520504731862,0.031545741324921134,0.21766561514195584,0.025236593059936908,0.0,0.12933753943217666,8,"['vlada.gov', 'www.faa.gov', 'www.cia.gov', 'www.cia.gov', 'webarchive.loc.gov', 'm.state.gov', 'www.cia.gov', 'www.cia.gov', 'uprava.gov', 'uprava.gov', 'www.britannica.com', 'www.bbc.com', 'economy.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.bbc.com', 'www.economist.com', 'books.google.com', 'www.euronews.com', 'www.nytimes.com', 'books.google.com', 'www.nytimes.com', 'www.pressreference.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'www.total-croatia-news.com', 'books.google.com', 'books.google.com', 'www.economist.com', 'www.aljazeera.com', 'www.nytimes.com', 'worldpopulationreview.com', 'articles.latimes.com', 'www.scribd.com', 'javno.com', 'books.google.com', 'www.nytimes.com', 'www.total-croatia-news.com', 'www.zgportal.com', 'articles.latimes.com', 'books.google.com', 'www.nytimes.com', 'www.nytimes.com', 'www.nytimes.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'setimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.styria.com', 'books.google.com', 'www.nytimes.com', 'www.nytimes.com', 'eurotestmobility.com', 'www.eubusiness.com', 'euro-poi.com', 'www.bbc.com', 'www.tehrantimes.com', 'books.google.com', 'www.total-croatia-news.com', 'www.nytimes.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'www.gallup.com', 'books.google.com', 'assets.pewresearch.org', 'www.eib.org', 'ourworldindata.org', 'go.worldbank.org', 'www.un.org', 'freedomhouse.org', 'whc.unesco.org', 'esa.un.org', 'ourworldindata.org', 'ourworldindata.org', 'h-net.org', 'ich.unesco.org', 'rsf.org', 'transparency.org', 'www.blueflag.org', 'www.un.org', 'jaspers.eib.org', 'datahelpdesk.worldbank.org', 'www.un.org', 'www.dubrovnik2011.sdewes.org', 'hdr.undp.org', 'milexdata.sipri.org', 'imf.org', ['bioscience'], ['unwto world tourism barometer '], ['european journal of international law'], ['revija za socijalnu politiku'], ['[[journal of genocide research'], ['acta medico-historica adriatica', 'hrvatsko znanstveno društvo za povijest zdravstvene kulture'], ['nature communications'], ['geoadria', 'hrvatsko geografsko društvo ']]",5573,Require administrator access (no expiry set),214161,3 September 2001,Koyaanis Qatsi ,11538,16,2001-09-03,2001-09,2001
180,180,Afghanistan,https://en.wikipedia.org/wiki/Afghanistan,521,10,"['10.3390/resources7030058', '10.1080/03068374.2015.1081001', '10.1038/s41467-020-19493-3', '10.1038/sdata.2018.214', '10.1371/journal.pone.0223111', '10.1080/07075332.1980.9640210', '10.1017/s1356186307007778', '10.1177/002200949703200207', '10.1007/s10680-005-6851-6', None, None, '33293507', '30375988', '31618275', None, None, None, None, None, None, '7723057', '6207062', '6795489', None, None, None, None]","[['resources'], ['asian affairs'], ['nature communications'], ['scientific data '], ['plos one'], ['the international history review '], ['journal of the royal asiatic society'], ['journal of contemporary history'], ['european journal of population']]",83,35,0,249,0,11,135,0.15930902111324377,0.0671785028790787,0.4779270633397313,0.019193857965451054,0.0,0.2456813819577735,9,"['pubs.usgs.gov', 'nato.usmission.gov', 'usaid.gov', 'pubs.usgs.gov', 'www.cia.gov', 'afghanistan.usaid.gov', 'afghanistan.usaid.gov', 'www.mfa.gov', 'prr.hec.gov', 'pubs.usgs.gov', '2009-2017.state.gov', 'pubs.usgs.gov', 'earthobservatory.nasa.gov', 'lcweb2.loc.gov', 'www.justice.gov', 'www.cia.gov', 'lcweb2.loc.gov', 'usaid.gov', 'webharvest.gov', 'www.mea.gov', 'pdf.usaid.gov', 'afghanistan.usaid.gov', 'www.mha.gov', 'pubs.usgs.gov', 'www.usaid.gov', 'www.cia.gov', 'prr.hec.gov', 'afghanistan.cr.usgs.gov', 'www.state.gov', 'www.dcda.gov', 'afghanistan.usaid.gov', 'pubs.usgs.gov', 'www.loc.gov', 'cia.gov', 'www.cia.gov', 'wadsam.com', 'www.news18.com', 'books.google.com', 'www.nytimes.com', 'www.afghanistans.com', 'messaging-custom-newsletters.nytimes.com', 'www.voanews.com', 'www.foxnews.com', 'www.thenation.com', 'www.afghan-web.com', 'ifpnews.com', 'designmena.com', 'www.nytimes.com', 'economictimes.indiatimes.com', 'statista.com', 'www.tolonews.com', 'www.bbc.com', 'news.yahoo.com', 'www.bbc.com', 'articles.latimes.com', 'thehill.com', 'www.tolonews.com', 'timesofindia.indiatimes.com', 'www.cbsnews.com', 'www.arabnews.com', 'edition.cnn.com', 'timesofindia.indiatimes.com', 'www.bt.com', 'www.bbc.com', 'encarta.msn.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.usatoday.com', 'www.pajhwok.com', 'www.afghan-web.com', 'www.aljazeera.com', 'books.google.com', 'www.cbsnews.com', 'books.google.com', 'www.youtube.com', 'www.reuters.com', 'www.dw.com', 'www.bloomberg.com', 'www.australiannationalreview.com', 'caravanistan.com', 'books.google.com', 'www.nytimes.com', 'amp.theaustralian.com', 'khorasanrugs.com', 'tribune.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.pajhwok.com', 'tribune.com', 'books.google.com', 'books.google.com', 'www.afghanistans.com', 'books.google.com', 'www.nytimes.com', 'www.cbsnews.com', 'www.nytimes.com', 'www.foodrepublic.com', 'www.afghanistans.com', 'tolonews.com', 'www.iexplore.com', 'books.google.com', 'www.aljazeera.com', 'www.papillonsartpalace.com', 'www.paulbogdanor.com', 'www.brecorder.com', 'www.afghanzariza.com', 'books.google.com', 'uk.reuters.com', 'tolonews.com', 'reference.com', 'edition.cnn.com', 'www.newstatesman.com', 'www.reuters.com', 'defenseindustrydaily.com', 'www.nytimes.com', 'www.dailyfinance.com', 'www.time.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.himalmag.com', 'books.google.com', 'en.mehrnews.com', 'www.britannica.com', 'www.nbcnews.com', 'infoplease.com', 'www.ft.com', 'www.dailytimes.com', 'bloomberg.com', 'reference.com', 'tolonews.com', 'www.cnbc.com', 'www.news18.com', 'ph.news.yahoo.com', 'www.youtube.com', 'bloomberg.com', 'www.nytimes.com', 'foreignpolicy.com', 'books.google.com', 'www.pajhwok.com', 'www.bbc.com', 'www.scmp.com', 'www.nytimes.com', 'books.google.com', 'books.google.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'ndtv.com', 'www.thehindu.com', 'books.google.com', 'www.britannica.com', 'www.reuters.com', 'www.redlandsdailyfacts.com', 'www.tolonews.com', 'referenceworks.brillonline.com', 'articles.chicagotribune.com', 'news.airwise.com', 'worldpopulationreview.com', 'thehill.com', 'www.reuters.com', 'www.hinduismtoday.com', 'www.nytimes.com', 'books.google.com', 'alamahabibi.com', 'www.voanews.com', 'www.aljazeera.com', 'www.bbc.com', 'www.teammelli.com', 'referenceworks.brillonline.com', 'books.google.com', 'www.youtube.com', 'www.csmonitor.com', 'books.google.com', 'worldpopulationreview.com', 'books.google.com', 'world.time.com', 'www.khaama.com', 'books.google.com', 'www.pajhwok.com', 'www.xinhuanet.com', 'www.msnbc.com', 'books.google.com', 'www.washingtonpost.com', 'www.wsj.com', 'www.nytimes.com', 'www.nytimes.com', 'articles.latimes.com', 'books.google.com', 'www.france24.com', 'books.google.com', 'www.nytimes.com', 'www.nytimes.com', 'books.google.com', 'www.telegraphindia.com', 'www.afghanistans.com', 'www.aljazeera.com', 'www.huffingtonpost.com', 'books.google.com', 'books.google.com', 'www.livemint.com', 'pajhwok.com', 'books.google.com', 'www.newsdaily.com', 'www.news18.com', 'books.google.com', 'books.google.com', 'bbcnazer.com', 'www.forbes.com', 'www.nytimes.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'www.csmonitor.com', 'books.google.com', 'tolonews.com', 'thediplomat.com', 'www.bbc.com', 'www.bbc.com', 'www.bbc.com', 'www.britannica.com', 'books.google.com', 'www.forbes.com', 'www.bbc.com', 'www.businessweek.com', 'www.afghanistans.com', 'afghan-web.com', 'www.bbc.com', 'books.google.com', 'www.washingtonpost.com', 'www.rareseeds.com', 'financialtribune.com', 'www.nytimes.com', 'books.google.com', 'www.voanews.com', 'www.bbc.com', 'www.soufangroup.com', 'books.google.com', 'news.yahoo.com', 'www.news24.com', 'edition.cnn.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.dw.com', 'tolonews.com', 'www.france24.com', 'www.csmonitor.com', 'books.google.com', 'measuredhs.com', 'www.bbc.com', 'www.bbc.com', 'www.economist.com', 'nl.newsbank.com', 'www.thehindu.com', 'www.topendsports.com', 'in.reuters.com', 'edition.cnn.com', 'acsor-surveys.com', 'thediplomat.com', 'books.google.com', 'www.france24.com', 'www.cnn.com', 'books.google.com', 'www.raillynews.com', 'bbcnazer.com', 'tolonews.com', 'www.trtworld.com', 'books.google.com', 'www.returntohope.com', 'www.raillynews.com', 'books.google.com', 'books.google.com', 'www.bangkokpost.com', 'afghanland.com', 'edition.cnn.com', 'books.google.com', 'www.brecorder.com', 'gandhara.com', 'abcnews.go.com', 'www.gounesco.com', 'daily.redbullmusicacademy.com', 'dictionary.cambridge.org', 'www.richardgregory.org', 'www.npr.org', 'www.pbs.org', 'nationalinterest.org', 'www.doctorswithoutborders.org', 'www.afghanistanjusticeproject.org', 'www.irinnews.org', 'www.asiafoundation.org', 'persian.packhum.org', 'gandhara.rferl.org', 'webarchive.urban.org', 'merip.org', 'www.unhcr.org', 'www.hrw.org', 'www.hrw.org', 'data.footprintnetwork.org', 'www.afghanistan-analysts.org', 'asiafoundation.org', 'news.un.org', 'www.rferl.org', 'www.afghanistan-analysts.org', 'philanthropynewsdigest.org', 'newsday.org', 'www.historycommons.org', 'data.worldbank.org', 'asiafoundation.org', 'persian.packhum.org', 'unama.unmissions.org', 'www.marxists.org', 'persian.packhum.org', 'www.afghanistan-analysts.org', 'seretandsons.org', 'www.irinnews.org', 'www.afghanistan-analysts.org', 'www.hrw.org', 'iranicaonline.org', 'www.imf.org', 'www.worldbank.org', 'www.medicamondiale.org', 'www.af.undp.org', 'www.prio.org', 'wayback.archive-it.org', 'en.unesco.org', 'www.prb.org', 'www.iranicaonline.org', 'wits.worldbank.org', 'www.afghanistanjusticeproject.org', 'data.worldbank.org', 'uis.unesco.org', 'monthlyreview.org', 'iec.org', 'www.hrw.org', 'www.npr.org', 'www.npr.org', 'www.nrfafg.org', 'freedomhouse.org', 'afghanistanembassy.org', 'globalvoices.org', 'www.pewforum.org', 'www.un.org', 'millenniumindicators.un.org', 'dictionary.cambridge.org', 'persian.packhum.org', 'www.rferl.org', 'data.worldbank.org', 'geonames.org', 'www.richardgregory.org', 'www.worldbank.org', 'www.afghanistan-analysts.org', 'publishing.cdlib.org', 'www.rferl.org', 'www.worldbank.org', 'www.unicef.org', 'uis.unesco.org', 'swedishcommittee.org', 'persian.packhum.org', 'hdr.undp.org', 'www.humandignitytrust.org', 'data.worldbank.org', 'www.afghanistan-analysts.org', 'publishing.cdlib.org', 'afghanistan.unfpa.org', ['resources'], ['asian affairs'], ['nature communications'], ['scientific data '], ['plos one'], ['the international history review '], ['journal of the royal asiatic society'], ['journal of contemporary history'], ['european journal of population']]",737,Require administrator access (no expiry set),297599,14 November 2001,Hagedis ,14819,34,2001-11-14,2001-11,2001
181,181,Sindhis,https://en.wikipedia.org/wiki/Sindhis,28,0,[],[],0,3,0,7,0,0,18,0.0,0.10714285714285714,0.25,0.0,0.0,0.10714285714285714,0,"['www.pbs.gov', 'www.censusindia.gov', 'lsi.gov', 'www.ethnologue.com', 'food.ndtv.com', 'www.newindianexpress.com', 'books.google.com', 'www.thenews.com', 'www.dawn.com', 'www.scribd.com']",446049,Allow all users (no expiry set),21909,28 January 2004,DigiBullet ,3997,9,2004-01-28,2004-01,2004
182,182,Poland,https://en.wikipedia.org/wiki/Poland,437,12,"['10.1017/s1014233900004582', '10.2307/3032734', '10.1080/00085006.1997.11092140', '10.1023/a:1007165901891', '10.1163/187633004x00116', '10.3917/poeu.021.0097', '10.1017/s0020818300006081', '10.1515/mgrsd-2017-0017', '10.14611/minib.21.09.2016.12', '10.1371/journal.pone.0054360', '10.1038/nature.2012.12020', '10.1080/0140238042000249876', None, None, None, None, None, None, None, None, None, '23342138', None, None, None, None, None, None, None, None, None, None, None, '3544712', None, None]","[['animal genetics resources information '], ['[[royal anthropological institute of great britain and ireland', '[[anthropology today'], ['[[taylor ', '[[canadian slavonic papers'], ['[[geojournal', '[[springer science'], [' east central europe '], ['politique européenne'], ['[[international organization ', '[[university of wisconsin press'], ['miscellanea geographica ', 'sciendo'], ['marketing of scientific and research organizations'], ['plos one '], ['nature news '], ['west european politics']]",44,38,0,198,0,3,142,0.10068649885583524,0.08695652173913043,0.45308924485125857,0.02745995423340961,0.0,0.2151029748283753,12,"['sejm.gov', 'stat.gov', 'aw.gov', 'stat.gov', 'isap.sejm.gov', 'www.cia.gov', 'stat.gov', 'stat.gov', 'psz.praca.gov', 'stat.gov', 'www.gov', 'www.paih.gov', 'gugik.gov', 'isap.sejm.gov', 'stat.gov', 'www.lasy.gov', 'www.stat.gov', 'www.parp.gov', 'stat.gov', 'ipn.gov', 'isap.sejm.gov', 'www.stat.gov', 'stat.gov', 'bip.cbsp.policja.gov', 'isap.sejm.gov', 'stat.gov', 'eteryt.stat.gov', 'www.gov', 'www.gddkia.gov', 'isap.sejm.gov', 'www.poland.gov', 'cba.gov', 'stat.gov', 'bip.mswia.gov', 'www.bbn.gov', 'orka.sejm.gov', 'isap.sejm.gov', 'www.mrr.gov', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.fifa.com', 'books.google.com', 'books.google.com', 'www.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.google.com', 'books.google.com', 'books.google.com', 'www.usnews.com', 'books.google.com', 'www.google.com', 'books.google.com', 'www.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.tourismroi.com', 'www.google.com', 'www.euromonitor.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thomaswhite.com', 'books.google.com', 'books.google.com', 'www.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.google.com', 'books.google.com', 'books.google.com', 'worldspeedway.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.xperiencepoland.com', 'geediting.com', 'www.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.slatkine.com', 'books.google.com', 'books.google.com', 'www.newgeography.com', 'www.google.com', 'www.google.com', 'emerging-europe.com', 'books.google.com', 'www.beautylish.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thoughtco.com', 'www.dw.com', 'www.expatica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.google.com', 'books.google.com', 'books.google.com', 'www.worldstopexports.com', 'books.google.com', 'www.dailysabah.com', 'www.google.com', 'italy-bulgaria2018.fivb.com', 'books.google.com', 'books.google.com', 'www.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.google.com', 'books.google.com', 'www.cnn.com', 'www.google.com', 'books.google.com', 'www.fifa.com', 'www.google.com', 'books.google.com', 'books.google.com', 'polandinexile.com', 'books.google.com', 'books.google.com', 'warsaw-life.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.google.com', 'books.google.com', 'justlanded.com', 'books.google.com', 'books.google.com', 'www.google.com', 'books.google.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'www.irishtimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.etymonline.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.etymonline.com', 'www.google.com', 'www.google.com', 'books.google.com', 'www.polandforvisitors.com', 'books.google.com', 'www.ft.com', 'www.google.com', 'books.google.com', 'books.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.janes.com', 'space.com', 'www.google.com', 'books.google.com', 'books.google.com', 'www.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.fivb.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.statista.com', 'www.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'countryeconomy.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.google.com', 'www.google.com', 'www.bbc.com', 'www.polishmeals.com', 'businessinsider.com', 'www.google.com', 'www.myjewishlearning.com', 'www.google.com', 'books.google.com', 'books.google.com', 'www.google.com', 'www.google.com', 'books.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.bbc.com', 'carnegieendowment.org', 'www.un.org', 'www.globalmethane.org', 'poland2014.fivb.org', 'data.worldbank.org', 'remember.org', 'stats.oecd.org', 'www.urbanaudit.org', 'hdr.undp.org', 'projectinposterum.org', 'www.sipri.org', 'siteresources.worldbank.org', 'read.oecd-ilibrary.org', 'www3.weforum.org', 'josephconradsociety.org', 'nobelprize.org', 'data.worldbank.org', 'encyclopedia.ushmm.org', 'www.gutenberg.org', 'npr.org', 'www.pisa.oecd.org', 'www.sat.org', 'encyclopedia.ushmm.org', 'data.worldbank.org', 'hdr.undp.org', 'www.yadvashem.org', 'whc.unesco.org', 'www2.unwto.org', 'data.worldbank.org', 'data.worldbank.org', 'data.worldbank.org', 'imf.org', 'rcin.org', 'data.worldbank.org', 'www.websters-online-dictionary.org', 'www.worldenergy.org', 'data.worldbank.org', 'josephconrad.org', 'hdr.undp.org', 'rynekpracy.org', 'www.oecd.org', 'data.worldbank.org', 'dataunodc.un.org', 'data.worldbank.org', ['animal genetics resources information '], ['[[royal anthropological institute of great britain and ireland', '[[anthropology today'], ['[[taylor ', '[[canadian slavonic papers'], ['[[geojournal', '[[springer science'], [' east central europe '], ['politique européenne'], ['[[international organization ', '[[university of wisconsin press'], ['miscellanea geographica ', 'sciendo'], ['marketing of scientific and research organizations'], ['plos one '], ['nature news '], ['west european politics']]",22936,Require administrator access (no expiry set),252203,13 November 2001,WojPob ,14351,50,2001-11-13,2001-11,2001
183,183,Georgia (country),https://en.wikipedia.org/wiki/Georgia_(country),350,4,"['10.1093/biosci/bix014', '10.1111/j.1468-2346.2008.00762.x', '10.1080/09668138808411783', '10.1038/s41467-020-19493-3', '28608869', None, None, '33293507', '5451287', None, None, '7723057']","[['bioscience'], ['[[international affairs '], ['soviet studies'], ['nature communications']]",72,29,0,61,0,3,181,0.2057142857142857,0.08285714285714285,0.1742857142857143,0.011428571428571429,0.0,0.3,4,"['government.gov', 'mfa.gov', 'mfa.gov', 'mod.gov', 'mfa.gov', 'tbilisi.gov', 'mreg.reestri.gov', 'mfa.gov', 'mfa.gov', 'mfa.gov', 'georgia.usembassy.gov', 'eia.doe.gov', 'www.president.gov', 'matsne.gov', 'mfa.gov', 'mes.gov', 'mfa.gov', 'www.smr.gov', 'www.loc.gov', 'delta.gov', 'matsne.gov', 'mfa.gov', 'www.cia.gov', 'mfa.gov', 'www.mes.gov', 'usa.mfa.gov', 'lcweb2.loc.gov', 'delta.gov', 'mfa.gov', 'www.bbc.com', 'foreignpolicy.com', 'rustavi2.com', 'topics.blogs.nytimes.com', 'books.google.com', 'www.reuters.com', 'books.google.com', 'www.washingtonpost.com', 'books.google.com', 'www.foxnews.com', 'www.rbth.com', 'books.google.com', 'www.forbes.com', 'www.bp.com', 'www.washingtonpost.com', 'www.rugbyworldcup.com', 'www.bbc.com', 'www.economist.com', 'books.google.com', 'rbedrosian.com', 'www.ft.com', 'www.bbc.com', 'search.ft.com', 'books.google.com', 'rbedrosian.com', 'www.britannica.com', 'www.reuters.com', 'www.reuters.com', 'books.google.com', 'cycloscope.weebly.com', 'edition.cnn.com', 'books.google.com', 'www.ukrferry.com', 'abcnews.go.com', 'online.wsj.com', 'search.ft.com', 'www.ukrferry.com', 'www.nytimes.com', 'www.britannica.com', 'www.euronews.com', 'www.bbc.com', 'findarticles.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'mcclatchydc.com', 'articles.chicagotribune.com', 'books.google.com', 'www.nytimes.com', 'www.bbc.com', 'www.hurriyetdailynews.com', 'www.bbc.com', 'newsru.com', 'ap.google.com', 'www.reuters.com', 'books.google.com', 'www.themoscowtimes.com', 'www.vinologue.com', 'www.ebrd.com', 'www.worldbank.org', 'hdr.undp.org', 'hdr.undp.org', 'www.rferl.org', 'www.rferl.org', 'cac-biodiversity.org', 'wayback.archive-it.org', 'eurasianet.org', 'wayback.archive-it.org', 'www.adb.org', 'imf.org', 'hrw.org', 'www.ndi.org', 'freedomhouse.org', 'www.unhcr.org', 'www.investingeorgia.org', 'www.eurasianet.org', 'data.worldbank.org', 'www.iri.org', 'wwf.panda.org', 'hrw.org', 'www.unesco.org', 'investingeorgia.org', 'data.worldbank.org', 'eurasianet.org', 'wayback.archive-it.org', 'www.leader.viitorul.org', 'www.crisisgroup.org', 'www.rferl.org', 'web.worldbank.org', 'www.pri.org', 'www.transparency.org', 'www.ge.undp.org', 'www.jamestown.org', 'www.rferl.org', 'jamestown.org', 'www.jamestown.org', 'wayback.archive-it.org', 'siteresources.worldbank.org', 'www.rferl.org', 'www.transparency.org', 'www.iucn.org', 'www.eurasianet.org', 'www.rferl.org', 'www.rferl.org', 'www.un.org', 'www.pirosmani.org', 'eurasianet.org', 'hrw.org', 'www.fidh.org', 'eurasianet.org', 'hrw.org', 'ich.unesco.org', 'www.doingbusiness.org', 'www.sss-tmas.org', 'www.worldbank.org', 'einung.org', 'ecmicaucasus.org', 'www.refworld.org', 'cybertruffle.org', 'hdr.undp.org', 'www.iranicaonline.org', 'cybertruffle.org', 'www.npr.org', 'freedomhouse.org', 'hrw.org', 'reports.weforum.org', 'www.napoleon-series.org', 'reports.weforum.org', 'osce.org', 'www.transparency.org', 'www.imf.org', ['bioscience'], ['[[international affairs '], ['soviet studies'], ['nature communications']]",48768,Require administrator access (no expiry set),225154,23 September 2001,Larry_Sanger ,10641,20,2001-09-23,2001-09,2001
184,184,Uzbekistan,https://en.wikipedia.org/wiki/Uzbekistan,256,5,"['10.1080/09662830008407454', '10.1086/342096', '10.1080/02634939608400946', '10.1093/biosci/bix014', '10.1093/jrs/4.4.372', None, '12145751', None, '28608869', None, None, '419996', None, '5451287', None]","[['european security'], ['the american journal of human genetics '], ['central asian survey '], ['bioscience'], ['journal of refugee studies ']]",77,14,0,72,0,5,84,0.30078125,0.0546875,0.28125,0.01953125,0.0,0.375,5,"['lcweb2.loc.gov', 'www.ustr.gov', 'www.cia.gov', 'usinfo.state.gov', 'data.gov', '2009-2017.state.gov', 'www.cia.gov', 'data.gov', 'data.gov', 'www.ustr.gov', 'data.gov', '2009-2017.state.gov', 'lcweb2.loc.gov', 'www.cia.gov', 'mecometer.com', 'www.thefreelibrary.com', 'www.cbsnews.com', 'www.nst.com', 'www.britannica.com', 'uzdaily.com', 'www.cbsnews.com', 'www.alamy.com', 'www.jweekly.com', 'www.business-anti-corruption.com', 'books.google.com', 'www.hsbc.com', 'www.orexca.com', 'www.the-afc.com', 'www.uzdaily.com', 'www.aljazeera.com', 'espn.com', 'uzwifi.com', 'www.bbc.com', 'enews.fergananews.com', 'books.google.com', 'www.c-and-a.com', 'www.newyorker.com', 'www.reuters.com', 'uzdaily.com', 'olympics.com', 'poltavareview.com', 'www.reuters.com', 'geopoliticalfutures.com', 'www.aljazeera.com', 'books.google.com', 'www.facebook.com', 'www.gazprom-international.com', 'www.uzdaily.com', 'www.eurasiareview.com', 'www.pilotguides.com', 'uzbek-travel.com', 'theglobaleconomy.com', 'www.cpamedia.com', 'bs-agro.com', 'books.google.com', 'www.globallegalinsights.com', 'chess.com', 'www.voanews.com', 'www.reuters.com', 'www.aa.com', 'www.bbc.com', 'www.voanews.com', 'worldatlas.com', 'factsanddetails.com', 'edition.cnn.com', 'www.chicagotribune.com', 'books.google.com', 'thediplomat.com', 'www.globallegalinsights.com', 'www.youtube.com', 'csrskabul.com', 'www.haaretz.com', 'cyclingtips.com', 'books.google.com', 'www.bbc.com', 'indexmundi.com', 'uzdaily.com', 'www.people-travels.com', 'www.newsweek.com', 'www.people-travels.com', 'time.com', 'www.forbes.com', 'www.time.com', 'www.teamuse.com', 'books.google.com', 'www.channelnewsasia.com', 'www.omct.org', 'www.rferl.org', 'data.worldbank.org', 'www.rferl.org', 'imf.org', 'www.world-nuclear.org', 'www.crisisgroup.org', 'hrw.org', 'tashkent.org', 'www.crisisgroup.org', 'databank.worldbank.org', 'eurasianet.org', 'www.rferl.org', 'www.ejfoundation.org', 'www.hrw.org', 'www.wilsoncenter.org', 'pewforum.org', 'www.aiba.org', 'www.doingbusiness.org', 'www.imf.org', 'eurasianet.org', 'bti-project.org', 'www.unhcr.org', 'web.amnesty.org', 'www.jewishvirtuallibrary.org', 'web.worldbank.org', 'investmentpolicyhub.unctad.org', 'www.cotton.org', 'globalslaveryindex.org', 'www.refworld.org', 'hdr.undp.org', 'www.globalpolicy.org', 'www.pewforum.org', 'news.trust.org', 'www.pewforum.org', 'www.the-sports.org', 'www.wto.org', 'www.amnesty.org', 'www.euronuclear.org', 'rsf.org', 'www.cacianalyst.org', 'voicesoncentralasia.org', 'data.worldbank.org', 'freedomhouse.org', 'www.rferl.org', 'www.imf.org', 'www.rferl.org', 'www.globalreligiousfutures.org', 'www.rferl.org', 'www.ihf-hr.org', 'www.osce.org', 'www.irinnews.org', 'hdr.undp.org', 'hdr.undp.org', 'www.msf.org', 'www.ihf-hr.org', 'kurash-ika.org', 'www.ajcarchives.org', 'www.rferl.org', 'www.aiba.org', 'uis.unesco.org', 'ilga.org', 'eurasiacenter.org', 'eurasianet.org', 'sdgs.un.org', 'collection.cooperhewitt.org', 'invest-in-uzbekistan.org', 'www.jamestown.org', 'adb.org', 'www.eurasianet.org', 'www.imf.org', 'kreml.org', 'www.iea.org', 'www.ajcarchives.org', 'rferl.org', 'www.ejfoundation.org', 'chalkboard.tol.org', ['european security'], ['the american journal of human genetics '], ['central asian survey '], ['bioscience'], ['journal of refugee studies ']]",31853,Require administrator access (no expiry set),161836,30 May 2001,KoyaanisQatsi ,7654,14,2001-05-30,2001-05,2001
185,185,Bosnia and Herzegovina,https://en.wikipedia.org/wiki/Bosnia_and_Herzegovina,230,4,"['10.1038/s41467-020-19493-3', '10.2307/3593383', '10.1093/biosci/bix014', '10.1075/lplp.28.1.03fai', '33293507', None, '28608869', None, '7723057', None, '5451287', None]","[['nature communications'], ['columbia law review', 'columbia law review association'], ['bioscience'], ['language problems ']]",29,8,0,81,0,3,105,0.12608695652173912,0.034782608695652174,0.3521739130434783,0.017391304347826087,0.0,0.1782608695652174,4,"['www.cia.gov', 'www.popis.gov', 'csce.gov', 'www.popis.gov', 'www.cia.gov', 'www.popis.gov', 'www.mod.gov', 'bhas.gov', 'books.google.com', 'books.google.com', 'public.dhe.ibm.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.globalfirepower.com', 'www.6yka.com', 'books.google.com', 'www.balkaninsight.com', 'books.google.com', 'encarta.msn.com', 'www.huffingtonpost.com', 'books.google.com', 'europeanwesternbalkans.com', 'apnews.com', 'ba.n1info.com', 'www.romereports.com', 'www.lonelyplanet.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.economist.com', 'books.google.com', 'www.tarasportrafting.com', 'books.google.com', 'www.aneks8komisija.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'ba.n1info.com', 'www.bbc.com', 'www.nezavisne.com', 'britannica.com', 'books.google.com', 'balkaninsight.com', 'books.google.com', 'www.reuters.com', 'getbybus.com', 'www.balkaninsight.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.smh.com', 'www.britannica.com', 'www.stripes.com', 'www.balkaninsight.com', 'features.us.reuters.com', 'www.internationalrafting.com', 'books.google.com', 'www.balkaninsight.com', 'reuters.com', 'ba.n1info.com', 'adventure.nationalgeographic.com', 'books.google.com', 'books.google.com', 'www.traveltalktours.com', 'books.google.com', 'books.google.com', 'books.google.com', 'courses.lumenlearning.com', 'foxnomad.com', 'www.scribd.com', 'books.google.com', 'www.britannica.com', 'www.economist.com', 'www.balkaninsight.com', 'businesswire.com', 'books.google.com', 'fuen.org', 'hdr.undp.org', 'data.worldbank.org', 'www.bosnia.org', 'iaaf.org', 'data.worldbank.org', 'data.worldbank.org', 'www.un.org', 'ufmsecretariat.org', 'hdr.undp.org', 'www.un.org', 'www.un.org', 'rsf.org', 'www.rferl.org', 'data.worldbank.org', 'www.ilo.org', 'un.org', 'phron.org', 'secnet069.un.org', 'www.hrw.org', 'www.un.org', 'www.rferl.org', 'www.un.org', 'www.pewforum.org', 'www.imf.org', 'rferl.org', 'hdr.undp.org', 'www.icty.org', 'ftp.fao.org', ['nature communications'], ['columbia law review', 'columbia law review association'], ['bioscience'], ['language problems ']]",3463,Require administrator access (no expiry set),208890,22 April 2001,Koyaanisqatsi ,10659,4,2001-04-22,2001-04,2001
186,186,Lebanon,https://en.wikipedia.org/wiki/Lebanon,365,7,"['10.1038/s41467-020-19493-3', '10.1177/001654928002600202', '10.1080/13642987.2017.1371140', '10.2307/2009820', '10.1093/jogss/ogz016', '10.1093/biosci/bix014', '10.1525/jps.1981.11.1.00p0366x', '33293507', None, None, None, None, '28608869', None, '7723057', None, None, None, None, '5451287', None]","[['nature communications'], ['gazette '], ['the international journal of human rights'], ['world politics'], ['journal of global security studies'], ['bioscience'], ['journal of palestine studies']]",63,35,0,151,0,1,109,0.1726027397260274,0.0958904109589041,0.4136986301369863,0.019178082191780823,0.0,0.2876712328767123,7,"['2001-2009.state.gov', '2009-2017.state.gov', 'www.lebarmy.gov', 'mfa.gov', 'www.cia.gov', 'www.lebanonundersiege.gov', 'www.lebarmy.gov', 'www.state.gov', 'www.cia.gov', '2009-2017.state.gov', 'www.moph.gov', 'www.cia.gov', 'www.moph.gov', 'webarchive.loc.gov', 'www.moph.gov', '2009-2017.state.gov', 'www.lebanon-tourism.gov', 'www.loc.gov', 'www.state.gov', 'www.fco.gov', '2009-2017.state.gov', 'hdl.loc.gov', 'lcweb2.loc.gov', 'hdl.loc.gov', 'www.mfa.gov', 'www.lebanonundersiege.gov', 'lebanon-tourism.gov', 'www.higher-edu.gov', 'export.gov', 'presidency.gov', 'destinationlebanon.gov', '2001-2009.state.gov', 'www.cia.gov', 'share.america.gov', 'www.cia.gov', 'www.aljazeera.com', 'books.google.com', 'www.bbc.com', 'www.nytimes.com', 'fiba.com', 'aljazeera.com', 'www.bbc.com', 'www.mtv.com', 'www.newyorker.com', 'about.com', 'www.time.com', 'www.hinduonnet.com', 'www.dailystar.com', 'www.dw.com', 'www.topuniversities.com', 'www.nationmaster.com', 'religionnews.com', 'www.washingtonpost.com', 'www.the961.com', 'www.france24.com', 'books.google.com', 'www.washingtonpost.com', 'www.dailystar.com', 'lebanonwaterfestival.com', 'www.dailystar.com', 'bbc.com', 'fanack.com', 'goalzz.com', 'www.dailystar.com', 'aljazeera.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.dailystar.com', 'apnews.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.dailystar.com', 'www.arabamerica.com', 'www.alyaum.com', 'www.thestar.com', 'abcnews.go.com', 'the961.com', 'www.ain-al-yaqeen.com', 'www.nytimes.com', 'thediplomat.com', 'books.google.com', 'yalla10.yalla.com', 'www.dailystar.com', 'www.reuters.com', 'voanews.com', 'www.dailystar.com', 'www.officeholidays.com', 'www.dailystar.com', 'www.dailystar.com', 'edition.cnn.com', 'www.reuters.com', 'www.newyorker.com', 'fanack.com', 'books.google.com', 'gulfnews.com', 'www.cynews.com', 'books.google.com', 'www.nytimes.com', 'www.smithsonianmag.com', 'www.cnn.com', 'www.dailystar.com', 'www.stratfor.com', 'www.dailystar.com', 'books.google.com', 'www.reuters.com', 'lebanonfiles.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'in.reuters.com', 'www.thenation.com', 'www.nytimes.com', 'www.al-monitor.com', 'www.iatatravelcentre.com', 'es.euronews.com', 'www.the961.com', 'www.topuniversities.com', 'www.opportunities.com', 'www.aljazeera.com', 'www.france24.com', 'www.naharnet.com', 'www.usatoday.com', 'books.google.com', 'books.google.com', 'www.time.com', 'www.dailystar.com', 'www.rsssf.com', 'www.aljazeera.com', 'www.britannica.com', 'www.idal.com', 'www.globalpolitician.com', 'en.mehrnews.com', 'kaftoun.com', 'football.com', 'books.google.com', 'books.google.com', 'bloomberg.com', 'dailystar.com', 'books.google.com', 'www.katagogi.com', 'www.nytimes.com', 'books.google.com', 'www.economist.com', 'fiba.com', 'www.rugbyleagueplanet.com', 'books.google.com', 'www.nytimes.com', 'www.audi.com', 'www.mtv.com', 'adcidl.com', 'www.deseretnews.com', 'www.dailystar.com', 'www.ehdenfamilytree.com', 'www.mallat.com', 'www.britannica.com', 'www.bbc.com', 'books.google.com', 'www.dailystar.com', 'articles.cnn.com', 'www.dailystar.com', 'fiba.com', 'bqdoha.com', 'www.the961.com', 'www.dailystar.com', 'lebanonwaterfestival.com', 'www.nytimes.com', 'www.couriermail.com', 'friesian.com', 'dailystar.com', 'www.france24.com', 'www.google.com', 'www.youtube.com', 'stepfeed.com', 'observers.france24.com', 'www.bbc.com', 'www.thenationalnews.com', 'www.topuniversities.com', 'www.middleeastmonitor.com', 'www.chron.com', 'www.the961.com', 'www.nytimes.com', 'books.google.com', 'abcnews.go.com', 'books.google.com', 'www.un.org', 'www.jta.org', 'domino.un.org', 'data2.unhcr.org', 'www.lstatic.org', 'www.hrw.org', 'www.usip.org', 'www.imf.org', 'www.un.org', 'data.worldbank.org', 'www.fao.org', 'www.hrw.org', 'data.worldbank.org', 'www.csbe.org', 'www.unesco.org', 'www.freedomhouse.org', 'www.hrw.org', 'www3.weforum.org', 'www.blueplanetbiomes.org', 'www.unhcr.org', 'www.tni.org', 'www.sesrtcic.org', 'stmaron.org', 'www.samidoun.org', 'carnegieendowment.org', 'www.usip.org', 'whc.unesco.org', 'www.amnesty.org', 'un.org', 'www.euroscience.org', 'beirutmarathon.org', 'www.rugbyleagueproject.org', 'www.irinnews.org', 'hrw.org', 'info.worldbank.org', 'www.cggl.org', 'data.worldbank.org', 'shoufcedar.org', 'www.carnegieendowment.org', 'www.evangelical-times.org', 'hdrstats.undp.org', 'www.npr.org', 'www.icrc.org', 'www.unhcr.org', 'www.irinnews.org', 'data.unhcr.org', 'www.libandata.org', 'www.pbs.org', 'www.carnegieendowment.org', 'www.worldvaluessurvey.org', 'www.pbs.org', 'www.olympic.org', 'nyulawglobal.org', 'www.sesrtcic.org', 'www.pogar.org', 'hdr.undp.org', 'www.jstor.org', 'www.un.org', 'washingtoninstitute.org', 'www.washingtoninstitute.org', 'www.pewresearch.org', 'www.foreignaffairs.org', 'un.org', ['nature communications'], ['gazette '], ['the international journal of human rights'], ['world politics'], ['journal of global security studies'], ['bioscience'], ['journal of palestine studies']]",17771,Allow all users (no expiry set),231802,18 May 2001,KoyaanisQatsi ,16844,14,2001-05-18,2001-05,2001
187,187,East India,https://en.wikipedia.org/wiki/East_India,97,0,[],[],6,16,0,54,0,0,21,0.061855670103092786,0.16494845360824742,0.5567010309278351,0.0,0.0,0.2268041237113402,0,"['tcpomud.gov', 'www.censusindia.gov', 'www.portal.gsi.gov', 'www.jharkhand.gov', 'census.gov', 'www.westbengaltourism.gov', 'tcpomud.gov', 'www.orissatourism.gov', 'www.westbengaltourism.gov', 'odishatourism.gov', 'southport.jpl.nasa.gov', 'orissa.gov', 'www.westbengal.gov', 'www.sundargarhzp.odishapr.gov', 'www.orissaminerals.gov', 'census.gov', 'www.telegraphindia.com', 'www.fifa.com', 'odissi.itgo.com', 'www.ccfc1792.com', 'books.google.com', 'articles.timesofindia.indiatimes.com', 'www.telegraphindia.com', 'm.bhaskar.com', 'www.indianexpress.com', 'books.google.com', 'www.nytimes.com', 'www.telegraphindia.com', 'www.hindu.com', 'books.google.com', 'www.fifa.com', 'www.hindu.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.aitatennis.com', 'www.hindustantimes.com', 'www.newindianexpress.com', 'orissalinks.com', 'www.telegraphindia.com', 'articles.timesofindia.indiatimes.com', 'in.news.yahoo.com', 'odishasuntimes.com', 'books.google.com', 'books.google.com', 'archive.wikiwix.com', 'rediff.com', 'www.telegraphindia.com', 'www.rugbyworldcup.com', 'books.google.com', 'books.google.com', 'articles.timesofindia.indiatimes.com', 'books.google.com', 'www.telegraphindia.com', 'books.google.com', 'thekalingalancers.com', 'timesofindia.indiatimes.com', 'www.telegraphindia.com', 'www.hindu.com', 'www.telegraphindia.com', 'www.espncricinfo.com', 'books.google.com', 'economictimes.indiatimes.com', 'books.google.com', 'theinfoindia.com', 'www.thehindu.com', 'dnaindia.com', 'www.hindustantimes.com', 'the-ifa.org', 'www.kmdaonline.org', 'www.metropolis.org', 'www.orissacricket.org', 'asiranchi.org', 'www.uraaei.org']",3799826,Allow all users (no expiry set),98982,21 January 2006,QuartierLatin1968 ,1663,5,2006-01-21,2006-01,2006
188,188,Belarus,https://en.wikipedia.org/wiki/Belarus,288,6,"['10.1108/978-1-83867-695-720191016', '10.1007/s12290-008-0029-7', '10.1080/1080/09668130500199509', '10.1093/biosci/bix014', '10.1080/15579336.2001.11770234', '10.1007/978-3-658-13762-5_19', None, None, None, '28608869', None, None, None, None, None, '5451287', None, None]","[['emerald publishing limited'], ['european view '], ['europe-asia studies '], ['bioscience'], ['international journal of sociology'], ['vergleichende politikwissenschaft. springer vs']]",39,35,0,94,0,2,112,0.13541666666666666,0.12152777777777778,0.3263888888888889,0.020833333333333332,0.0,0.2777777777777778,6,"['cia.gov', 'www.mfa.gov', 'mfa.gov', 'www.cia.gov', 'belstat.gov', 'www.cia.gov', 'www.cia.gov', 'president.gov', 'usinfo.state.gov', 'census.belstat.gov', 'mfa.gov', 'www.president.gov', 'president.gov', 'www.cia.gov', 'www.belstat.gov', 'www.minsk.gov', 'www.cia.gov', 'www.census.gov', 'www.gov', 'www.belstat.gov', 'www.belstat.gov', 'belstat.gov', 'www.president.gov', 'rec.gov', 'www.mfa.gov', 'president.gov', '2009-2017.state.gov', 'www.president.gov', 'www.mrik.gov', '2009-2017.state.gov', 'english.gov', 'www.mfa.gov', 'mfa.gov', 'www.minsk.gov', 'president.gov', 'foreignpolicy.com', 'www.worldatlas.com', 'books.google.com', 'www.business-anti-corruption.com', 'fotw.fivestarflags.com', 'www.voanews.com', 'www.reuters.com', 'books.google.com', 'www.msn.com', 'books.google.com', 'www.belarusguide.com', 'www.nationmaster.com', 'www.wsj.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'belarus-travel.com', 'belarusguide.com', 'www.reuters.com', 'world-gazetteer.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'www.themoscowtimes.com', 'www.statista.com', 'www.stalbertgazette.com', 'www.nationmaster.com', 'www.smh.com', 'www.nytimes.com', 'app1.chinadaily.com', 'www.nytimes.com', 'books.google.com', 'www.nbcnews.com', 'books.google.com', 'apnews.com', 'www.voiceofbelarus.com', 'www.books-by-isbn.com', 'www.kyivpost.com', 'books.google.com', 'www.bbc.com', 'books.google.com', 'www.euronews.com', 'www.nytimes.com', 'www.reuters.com', 'books.google.com', 'books.google.com', 'apnews.com', 'belarusguide.com', 'books.google.com', 'www.vice.com', 'ethnologue.com', 'books.google.com', 'www.dw.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'pravo.kulichki.com', 'books.google.com', 'www.dw.com', 'books.google.com', 'books.google.com', 'news.sky.com', 'books.google.com', 'books.google.com', 'uk.reuters.com', 'books.google.com', 'books.google.com', 'euobserver.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.washingtonpost.com', 'www.axios.com', 'news.yahoo.com', 'france24.com', 'www.euronews.com', 'www.ft.com', 'foreignpolicy.com', 'books.google.com', 'landofancestors.com', 'content.time.com', 'notesfrompoland.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'books.google.com', 'seattletimes.com', 'www.nytimes.com', 'books.google.com', 'www.yahoo.com', 'timeanddate.com', 'books.google.com', 'books.google.com', 'britannica.com', 'chernobyl.undp.org', 'rferl.org', 'adsdatabase.ohchr.org', 'www.orfonline.org', 'charter97.org', 'wto.org', 'www.un.org', 'www.belarusembassy.org', 'hrw.org', 'jamestown.org', 'www.olympic.org', 'www.constituteproject.org', 'rsf.org', 'www.atlanticcouncil.org', 'www.osce.org', 'www.imf.org', 'tc.iaea.org', 'yivoencyclopedia.org', 'nobelprize.org', 'hrw.org', 'www.amnesty.org', 'www.fao.org', 'hdr.undp.org', 'www.un.org', 'www.amnesty.org', 'www.rferl.org', 'whc.unesco.org', 'currency-iso.org', 'www.heritage.org', 'hdr.undp.org', 'www.hrw.org', 'www.ohchr.org', 'data.worldbank.org', 'lnweb18.worldbank.org', 'www.rferl.org', 'data.worldbank.org', 'www.un.org', 'ru.forsecurity.org', 'kamunikat.org', ['emerald publishing limited'], ['european view '], ['europe-asia studies '], ['bioscience'], ['international journal of sociology'], ['vergleichende politikwissenschaft. springer vs']]",3457,Require autoconfirmed or confirmed access (no expiry set),162964,18 August 2001,Taw ,7797,7,2001-08-18,2001-08,2001
189,189,Aurangabad,https://en.wikipedia.org/wiki/Aurangabad,67,4,"['10.1017/cbo9780511576867.009', '10.4324/9780203483282-9', '10.1093/acprof:oso/9780190222536.001.0001', '10.1093/acprof:oso/9780190222536.003.0005', None, None, None, None, None, None, None, None]","[['cambridge university press'], ['routledge'], ['oxford university press'], ['oxford university press']]",7,13,0,16,0,0,27,0.1044776119402985,0.19402985074626866,0.23880597014925373,0.05970149253731343,0.0,0.3582089552238806,4,"['www.maharashtra.gov', 'censusindia.gov', 'census.gov', 'aurangabadcitypolice.gov', 'www.censusindia.gov', 'aurangabad.nielit.gov', 'aurangabad.gov', 'imdpune.gov', 'censusindia.gov', 'aurangabad.gov', 'imdpune.gov', 'aurangabad.gov', 'www.maharashtra.gov', 'economictimes.indiatimes.com', 'timesofindia.indiatimes.com', 'www.aurangabaddirectory.com', 'www.deccanherald.com', 'maharashtratimes.indiatimes.com', 'timesofindia.indiatimes.com', 'bangalorenotes.com', 'books.google.com', 'www.dnaindia.com', 'articles.timesofindia.indiatimes.com', 'economictimes.indiatimes.com', 'timesofindia.indiatimes.com', 'www.britannica.com', 'www.asianage.com', 'www.uppercrustindia.com', 'www.lokmat.com', 'jamaat.org', 'www.worldcat.org', 'www.cbaurangabad.org', 'www.worldcat.org', 'www.worldcat.org', 'jamaat.org', 'worldcat.org', ['cambridge university press'], ['routledge'], ['oxford university press'], ['oxford university press']]",546024,Allow all users (no expiry set),55631,23 March 2004,Hemanshu ,4645,14,2004-03-23,2004-03,2004
190,190,Azerbaijan,https://en.wikipedia.org/wiki/Azerbaijan,382,10,"['10.1093/biosci/bix014', '10.1017/s0041977x00090182', '10.1017/s0020743800064473', '10.3390/resources7030058', '10.1177/002200940103600202', '10.1038/s41467-020-19493-3', '10.1080/00210862.2020.1865136', '10.1038/sdata.2018.214', '10.1016/j.postcomstud.2013.09.001', '10.1057/978-1-137-38781-3_4', '28608869', None, None, None, None, '33293507', None, '30375988', None, None, '5451287', None, None, None, None, '7723057', None, '6207062', None, None]","[['bioscience'], ['bulletin of the school of oriental and african studies'], ['international journal of middle east studies'], ['resources'], ['journal of contemporary history '], ['nature communications'], ['iranian studies '], ['scientific data '], ['communist and post-communist studies '], ['[[palgrave macmillan']]",93,25,0,103,0,2,152,0.24345549738219896,0.06544502617801047,0.2696335078534031,0.02617801047120419,0.0,0.33507853403141363,10,"['www.loc.gov', 'stat.gov', 'www.fco.gov', '2017.state.gov', 'evisa.gov', 'baku.mfa.gov', 'www.mfa.gov', 'www.cia.gov', 'state.gov', 'www.dol.gov', 'www.diaspora.gov', 'www.loc.gov', 'cia.gov', 'ntrc.gov', 'courts.gov', 'www.mfa.gov', 'www.cia.gov', 'www.meclis.gov', 'lcweb2.loc.gov', 'www.stat.gov', 'cia.gov', 'www.dtxk.gov', 'www.cia.gov', 'www.cia.gov', 'www.state.gov', 'apnews.com', 'books.google.com', 'arthistoryarchive.com', 'www.ethnologue.com', 'books.google.com', 'azer.com', 'www.washingtonpost.com', 'www.google.com', 'www.britannica.com', 'www.bp.com', 'www.breakingisraelnews.com', 'www.nationsencyclopedia.com', 'www.hurriyetdailynews.com', 'www.vomcanada.com', 'www.azhydromet.com', 'baku2015.com', 'www.uefa.com', 'books.google.com', 'www1.chinadaily.com', 'www.reuters.com', 'books.google.com', 'edition.cnn.com', 'irs-az.com', 'www.space-travel.com', 'books.google.com', 'www.economist.com', 'www.dw.com', 'reports.chessdom.com', 'www.bbc.com', 'www.washingtontimes.com', 'encyclopedia2.thefreedictionary.com', 'worldatlas.com', 'www.google.com', 'www.satellitetoday.com', 'books.google.com', 'www.britannica.com', 'euobserver.com', 'azer.com', 'books.google.com', 'www.gallup.com', 'books.google.com', 'azer.com', 'www.uefa.com', 'worldatlas.com', 'www.azembassy.com', 'azer.com', 'books.google.com', 'brittanica.com', 'books.google.com', 'azer.com', 'www.britannica.com', 'www.nationsencyclopedia.com', 'books.google.com', 'www.keesings.com', 'www.theweekinchess.com', 'bp.com', 'books.google.com', 'www.forbes.com', 'www.window2baku.com', 'www.hurriyetdailynews.com', 'books.google.com', 'www.baku2017.com', 'books.google.com', 'books.google.com', 'books.google.com', 'apnews.com', 'books.google.com', 'www.bp.com', 'www.prweb.com', 'books.google.com', 'ru.uefa.com', 'www.fifa.com', 'books.google.com', 'nl.newsbank.com', 'www.thenationalnews.com', 'books.google.com', 'books.google.com', 'foreignpolicy.com', 'www.nytimes.com', 'en.clubatleticodemadrid.com', '(www.dw.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.washingtonpost.com', 'azer.com', 'books.google.com', 'www.dw.com', 'www.britannica.com', 'books.google.com', 'www.constructiondigital.com', 'books.google.com', 'www.time.com', 'books.google.com', 'books.google.com', 'www.com', 'www.azer.com', 'pqasb.pqarchiver.com', 'books.google.com', 'select.nytimes.com', 'www.newsweek.com', 'karabakhfoundation.org', 'www.catholic-hierarchy.org', 'rsf.org', 'www.azadliq.org', 'seismonet.org', 'fivb.org', 'www.azstat.org', 'data.un.org', 'www.amnesty.org', 'jns.org', 'www.iranicaonline.org', 'www.globalsocialscience.org', 'www.azstat.org', 'www.iranicaonline.org', 'www.doingbusiness.org', 'www.iranicaonline.org', 'www.eurasianet.org', 'passportindex.org', 'www.avesta.org', 'www.worldbank.org', 'www.un-az.org', 'www.rferl.org', 'www.un.org', 'cpj.org', 'www.worldbank.org', 'eurasianet.org', 'portal.unesco.org', 'www.iranicaonline.org', 'www.silkroadstudies.org', 'old.freedomhouse.org', 'www.keston.org', 'old.freedomhouse.org', 'www.cfom.org', 'www.doingbusiness.org', 'hdr.undp.org', 'hrw.org', 'imf.org', 'www.un.org', 'www.un.org', 'www.eurolympic.org', 'www.hrw.org', 'www.esiweb.org', 'azstat.org', 'unstats.un.org', 'www.eurasianet.org', 'www.hrw.org', 'nkrusa.org', 'www.osce.org', 'www3.weforum.org', 'peacemaker.un.org', 'www.hrw.org', 'data.footprintnetwork.org', 'universes-in-universe.org', 'features.pewforum.org', 'www.silkroadstudies.org', 'azstat.org', 'peacemaker.un.org', 'www.rferl.org', 'pewforum.org', 'www.amnesty.org', 'esisc.org', 'whc.unesco.org', 'freedomhouse.org', 'www.azstat.org', 'library.aliyev-heritage.org', 'www.jta.org', 'pewforum.org', 'www.unesco.org', 'wttc.org', 'www.un.org', 'worldheritagesite.org', 'www.eurasianet.org', 'www.cac-biodiversity.org', 'www.freedomhouse.org', 'www.refworld.org', 'www3.weforum.org', 'freedomhouse.org', 'www.un.org', 'esisc.org', 'www.un-az.org', 'www.worldheritagesite.org', 'www.eurasianet.org', 'ask.org', 'eanpages.org', 'www.azstat.org', 'www.silkroadstudies.org', 'www.jewishvirtuallibrary.org', 'www.eurasianet.org', 'civicsolidarity.org', 'hdr.undp.org', 'www.un.org', 'www.cac-biodiversity.org', 'www.jamestown.org', ['bioscience'], ['bulletin of the school of oriental and african studies'], ['international journal of middle east studies'], ['resources'], ['journal of contemporary history '], ['nature communications'], ['iranian studies '], ['scientific data '], ['communist and post-communist studies '], ['[[palgrave macmillan']]",746,Require administrator access (no expiry set),237548,31 October 2001,Corvus13 ,10120,22,2001-10-31,2001-10,2001
191,191,Amatrice,https://en.wikipedia.org/wiki/Amatrice,9,0,[],[],0,0,0,4,0,1,4,0.0,0.0,0.4444444444444444,0.0,0.0,0.0,0,"['www.reuters.com', 'edition.cnn.com', 'www.portaleabruzzo.com', 'www.bbc.com']",5710172,Allow all users (no expiry set),11205,25 June 2006,Attilios ,271,0,2006-06-25,2006-06,2006
192,192,Chumash people,https://en.wikipedia.org/wiki/Chumash_people,92,9,"['10.1007/bf00889174', '10.1007/bf02860489', '10.1093/ecam/nem188', '10.2307/40035309', '10.1093/ecam/neh090', '10.2307/2694568', '10.1525/aa.2005.107.3.432', '10.1353/aiq.2006.0020', '10.1525/aa.1995.97.4.02a00150', None, None, '18955312', None, '15937554', None, None, None, None, None, None, '2862936', None, '1142202', None, None, None, None]","[[' human ecology '], [' [[economic botany'], ['evidence-based complementary and alternative medicine'], ['american antiquity'], [' evidence-based complementary and alternative medicine'], [' american antiquity '], ['american anthropologist', 'american anthropological association'], [' american indian quarterly '], [' american anthropologist ']]",11,7,0,14,0,0,51,0.11956521739130435,0.07608695652173914,0.15217391304347827,0.09782608695652174,0.0,0.29347826086956524,9,"['www.nps.gov', 'ftp.consrv.ca.gov', 'www.nps.gov', 'www.loc.gov', 'www.nps.gov', 'ftp.consrv.ca.gov', 'www.nps.gov', 'www.reuters.com', 'content.time.com', 'books.google.com', 'sanluisobispo.com', 'www.latimes.com', 'www.nwmarinelife.com', 'www.mercurynews.com', 'www.sfgate.com', 'wildfoodplants.com', 'donnamiscolta.com', 'ranchopalosverdes.patch.com', 'www.youtube.com', 'www.independent.com', 'sanluisobispo.com', 'www.wishtoyo.org', 'calisphere.org', 'www.santaynezchumash.org', 'syceo.org', 'americanindian2.abc-clio.com.libaccess.sjlibrary.org', 'www.pcas.org', 'www.seathos.org', 'calisphere.org', 'www.wishtoyo.org', 'www.veggierescue.org', 'www.sbnature.org', [' human ecology '], [' [[economic botany'], ['evidence-based complementary and alternative medicine'], ['american antiquity'], [' evidence-based complementary and alternative medicine'], [' american antiquity '], ['american anthropologist', 'american anthropological association'], [' american indian quarterly '], [' american anthropologist ']]",92492,Allow all users (no expiry set),62051,26 September 2002,David depaoli ,1409,10,2002-09-26,2002-09,2002
193,193,Culture of Armenia,https://en.wikipedia.org/wiki/Culture_of_Armenia,17,0,[],[],1,1,0,6,0,0,9,0.058823529411764705,0.058823529411764705,0.35294117647058826,0.0,0.0,0.11764705882352941,0,"['www.gov', 'www.imdb.com', 'www.egofilmarts.com', 'www.nayiri.com', 'bayrakdarian.com', 'www.armenmusic.com', 'armeniansongbook.com', 'www.unesco.org']",2049464,Allow all users (no expiry set),25973,15 June 2005,Protarion ,676,1,2005-06-15,2005-06,2005
194,194,Huế,https://en.wikipedia.org/wiki/Hu%E1%BA%BF,44,0,[],[],5,0,0,7,0,0,32,0.11363636363636363,0.0,0.1590909090909091,0.0,0.0,0.11363636363636363,0,"['www.huesmiletravel.com', 'travel-tourist-information-guide.com', 'asiamarvels.com', 'www.bangkokbiznews.com', 'www.gonomad.com', 'www.thingsasian.com', 'www.aftabir.com', 'plumvillage.org', 'whc.unesco.org', 'www.sister-cities.org', 'cdkn.org', 'cdkn.org']",59684,Allow all users (no expiry set),41617,27 June 2002,203.109.250.99 ,1204,3,2002-06-27,2002-06,2002
195,195,Armenia,https://en.wikipedia.org/wiki/Armenia,249,5,"['10.3390/resources7030058', '10.5281/zenodo.1240524', '10.1093/acref/9780199546091.001.0001', '10.1093/biosci/bix014', '10.1038/sdata.2018.214', None, None, None, '28608869', '30375988', None, None, None, '5451287', '6207062']","[['resources '], ['zenodo '], ['[[cia', '[[national geographic society', 'istituto geografico de agostini', 'oxford reference online '], ['bioscience'], ['scientific data ']]",36,12,0,59,0,1,137,0.14457831325301204,0.04819277108433735,0.23694779116465864,0.020080321285140562,0.0,0.21285140562248997,5,"['www.mfa.gov', 'www.mfa.gov', 'www.cia.gov', 'webarchive.loc.gov', 'www.census.gov', 'cia.gov', 'lcweb2.loc.gov', 'www.cia.gov', 'www.cia.gov', 'www.gov', 'www.gov', 'www.census.gov', 'books.google.com', 'www.bolsohays.com', 'www.todayszaman.com', 'books.google.com', 'www.smithsonianmag.com', 'dictionary.com', 'news.nationalgeographic.com', 'www.goodnewsadvertising.com', 'apnews.com', 'books.google.com', 'www.google.com', 'www.google.com', 'www.countriesquest.com', 'cdn.discordapp.com', 'www.theglobeandmail.com', 'www.dw.com', 'books.google.com', 'ancienthistory.about.com', 'europeforvisitors.com', 'books.google.com', 'books.google.com', 'www.aljazeera.com', 'www.britannica.com', 'books.google.com', 'gallup.com', 'books.google.com', 'books.google.com', 'books.google.com', 'farm1.staticflickr.com', 'www.nationalgeographic.com', 'www.pseudepigrapha.com', 'www.newindianexpress.com', 'news.yahoo.com', 'books.google.com', 'www.aljazeera.com', 'books.google.com', 'www.armenianow.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.cnn.com', 'encyclopedia2.thefreedictionary.com', 'www.economist.com', 'www.aljazeera.com', 'www.libertas-institut.com', 'www.google.com', 'www.washingtonpost.com', 'www.aa.com', 'books.google.com', 'www.highbeam.com', 'books.google.com', 'welcomearmenia.com', 'www.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.worldhistory.org', 'data.footprintnetwork.org', 'aceproject.org', 'www.globalheritagefund.org', 'fragilestatesindex.org', 'www.fraserinstitute.org', 'www.minorities-network.org', 'freedomhouse.org', 'www.armenian-genocide.org', 'www.soviethistory.org', 'unesdoc.unesco.org', 'imf.org', 'hdr.undp.org', 'www.crisisgroup.org', 'www.rferl.org', 'rsf.org', 'rsf.org', 'abcy.org', 'www.cato.org', 'rsf.org', 'www.rferl.org', 'www.eurasianet.org', 'www.jewishvirtuallibrary.org', 'visitarmenia.org', 'cato.org', 'hdr.undp.org', 'www.eurasiancommission.org', 'freedomhouse.org', 'www.constituteproject.org', 'www.rferl.org', 'data.worldbank.org', 'fragilestatesindex.org', 'www.heritage.org', 'rsf.org', 'www.armenianchurch.org', 'www.cfr.org', ['resources '], ['zenodo '], ['[[cia', '[[national geographic society', 'istituto geografico de agostini', 'oxford reference online '], ['bioscience'], ['scientific data ']]",10918072,Require administrator access (no expiry set),192345,2 July 2001,KoyaanisQatsi ,7924,13,2001-07-02,2001-07,2001
196,196,Coastal Andhra,https://en.wikipedia.org/wiki/Coastal_Andhra,15,0,[],[],0,3,0,9,0,0,3,0.0,0.2,0.6,0.0,0.0,0.2,0,"['dof.gov', 'www.ap.gov', 'censusindia.gov', 'www.thehindu.com', 'www.preservearticles.com', 'www.livemint.com', 'mapsofindia.com', 'www.mapsofindia.com', 'www.business-standard.com', 'www.thehindu.com', 'books.google.com', 'www.thehindu.com']",990249,Allow all users (no expiry set),18111,16 September 2004,Tom Radulovich ,931,7,2004-09-16,2004-09,2004
197,197,Bologna,https://en.wikipedia.org/wiki/Bologna,116,0,[],[],7,2,0,22,0,0,86,0.0603448275862069,0.017241379310344827,0.1896551724137931,0.0,0.0,0.07758620689655173,0,"['2001-2009.state.gov', 'www.gov', 'books.google.com', 'www.metro-report.com', 'www.experiencefestival.com', 'www.baseballprospectus.com', 'www.topuniversities.com', 'www.ilsole24ore.com', 'www.espn.com', 'books.google.com', 'cittadellamusica.com', 'moovitapp.com', 'artcityemiliaromagna.com', 'aaa-angelica.com', 'www.unicreditreviews.com', 'www.com', 'www.com', 'www.fortitudobaseball.com', 'www.unicreditreviews.com', 'www.citymayors.com', 'www.someprefercakefestival.com', 'books.google.com', 'books.google.com', 'moovitapp.com', 'whc.unesco.org', 'portal.unesco.org', 'climaintoscana.altervista.org', 'futurefilmfestival.org', 'www.yesmagazine.org', 'www.italo-americana.org', 'creativecommons.org']",21069333,Allow all users (no expiry set),94523,25 February 2002,MichaelTinkler ,3152,7,2002-02-25,2002-02,2002
198,198,Romani people,https://en.wikipedia.org/wiki/Romani_people,302,20,"['10.1002/ajpa.21372', '10.1086/324681', '10.1017/s2071832200005423', '10.1093/molbev/msi185', '10.15196/ts580101', '10.3389/fgene.2019.00558', '10.1038/sj.ejhg.5200597', '10.1371/journal.pone.0048477', '10.1038/ejhg.2015.201', '10.1186/1471-2350-2-5', '10.1093/molbev/msaa156', '10.1016/j.cub.2012.10.039', '10.1537/ase.090203', None, '10.1371/journal.pone.0056779', '10.1086/424759', '10.1111/j.1469-1809.2005.00251.x', '10.1016/j.fsigen.2014.06.013', '10.1080/0032472031000147856', '10.1038/nature02029', '20878647', '11704928', None, '15944443', None, '31263480', '11313742', '23209554', '26374132', '11299048', '32589725', '23219723', None, None, '23483890', '15322984', '16759179', '25051224', None, '14647380', None, '1235543', None, None, None, '6585392', None, '3509117', '4867443', '31389', None, None, None, 'year', '3590186', '1182047', None, '4234079', None, None]","[['american journal of physical anthropology '], [' american journal of human genetics '], ['german law journal '], [' mol. biol. evol. '], [' területi statisztika '], ['frontiers in genetics '], ['european journal of human genetics '], [' plos one '], ['european journal of human genetics '], ['bmc medical genetics '], ['molecular biology and evolution'], ['current biology '], ['anthropological science '], [' univ of hertfordshire press '], [' plos one '], ['the american journal of human genetics '], ['annals of human genetics '], [' forensic science international. genetics '], [' population studies '], [' [[nature ']]",37,9,0,72,0,4,161,0.12251655629139073,0.029801324503311258,0.23841059602649006,0.06622516556291391,0.0,0.2185430463576159,20,"['www.stat.gov', 'belstat.gov', 'webrzs.stat.gov', 'dane.gov', 'www.nyed.uscourts.gov', '2001.ukrcensus.gov', 'www.america.gov', 'instat.gov', 'www.msd.gov', 'www.ethnologue.com', 'www.iranian.com', 'books.google.com', 'theconversation.com', 'www.isidore-of-seville.com', 'india.com', 'www.reuters.com', 'www.scritub.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'kopachi.com', 'www.dw.com', 'www.etymonline.com', 'hindugateway.com', 'www.euractiv.com', 'books.google.com', 'www.thefreedictionary.com', 'www.aljazeera.com', 'books.google.com', 'greece.greekreporter.com', 'www.geocities.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'eupedia.com', 'books.google.com', 'www.geocities.com', 'books.google.com', 'www.livescience.com', 'www.wernercohn.com', 'apnews.com', 'books.google.com', 'books.google.com', 'www.csmonitor.com', 'www.nytimes.com', 'elpais.com', 'usatoday30.usatoday.com', 'www.youscribe.com', 'books.google.com', 'books.google.com', 'www.everyculture.com', 'books.google.com', 'webarsiv.hurriyet.com', 'www.rootsworld.com', 'www.reocities.com', 'www.omniglot.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.milliyet.com', 'books.google.com', 'books.google.com', 'www.khaleejtimes.com', 'www.everyculture.com', 'www.ethnologue.com', 'books.google.com', 'noticias.r7.com', 'english.elpais.com', 'www.heyalma.com', 'www.tlc.com', 'content.time.com', 'books.google.com', 'www.nytimes.com', 'usatoday30.usatoday.com', 'books.google.com', 'www.la-croix.com', 'www.ethnologue.com', 'books.google.com', 'draganprimorac.com', 'www.bbc.com', 'www.undv.org', 'www.florilegium.org', 'www.eumap.org', 'www.ushmm.org', 'www.monstat.org', 'www.iranicaonline.org', 'journals.plos.org', 'www.restlessbeings.org', 'www.gypsyloresociety.org', 'opensourcefoundations.org', 'minorityrights.org', 'www.balkanproject.org', 'www.pewresearch.org', 'www.wiseattention.org', 'www.amnesty.org', 'www.oikoumene.org', 'newsdesk.org', 'www.refworld.org', 'www.21luglio.org', 'web.amnesty.org', 'desicritics.org', 'theyliewedie.org', 'www.ushmm.org', 'www.errc.org', 'www.unhcr.org', 'www.pewglobal.org', 'romania.europalibera.org', 'www.rferl.org', 'holocaustcenter.jfcs.org', 'www.iranicaonline.org', 'www.radionetherlandsarchives.org', 'dhnet.org', 'www.berlin-institut.org', 'www.sca.org', 'www.errc.org', 'web.worldbank.org', 'www.savior.org', ['american journal of physical anthropology '], [' american journal of human genetics '], ['german law journal '], [' mol. biol. evol. '], [' területi statisztika '], ['frontiers in genetics '], ['european journal of human genetics '], [' plos one '], ['european journal of human genetics '], ['bmc medical genetics '], ['molecular biology and evolution'], ['current biology '], ['anthropological science '], [' univ of hertfordshire press '], [' plos one '], ['the american journal of human genetics '], ['annals of human genetics '], [' forensic science international. genetics '], [' population studies '], [' [[nature ']]",26152,Require administrator access (no expiry set),190289,15 November 2001,65.68.87.xxx ,10489,36,2001-11-15,2001-11,2001
199,199,Rome,https://en.wikipedia.org/wiki/Rome,198,6,"['10.1017/s0009840x00221331', '10.1177/1474885107080651', '10.2307/295257', '10.1086/361701', '10.1111/j.1468-2427.2010.00993.x', '10.1017/s0003598x00085859', None, None, None, None, None, None, None, None, None, None, None, None]","[['the classical review '], ['european journal of political theory '], ['the american journal of philology '], ['classical philology ', 'university of chicago press '], ['international journal of urban and regional research '], ['antiquity ', 'cambridge university press ']]",27,5,0,51,0,4,107,0.13636363636363635,0.025252525252525252,0.25757575757575757,0.030303030303030304,0.0,0.1919191919191919,6,"['www.tirana.gov', 'www.nyc.gov', 'www.ebeijing.gov', 'www.commune-tunis.gov', 'www.tirana.gov', 'www.britannica.com', 'www.mandatory.com', 'www.com', 'fendi.com', 'books.google.com', 'www.com', 'media.johnwiley.com', 'www.com', 'archive.wikiwix.com', 'initaly.com', 'www.washingtonpost.com', 'www.kurdishquestion.com', 'books.google.com', 'www.forbes.com', 'maspostatevilaregina.com', 'eurostar-av.trenitalia.com', 'www.romefile.com', 'www.questia.com', 'www.nytimes.com', 'www.cnn.com', 'guinnesworldrecords.com', 'www.com', 'www.historytoday.com', 'languagemonitor.com', 'www.com', 'www.visiterome.com', 'www.ilsole24ore.com', 'www.com', 'www.citymayors.com', 'www.rometales.com', 'history.com', 'www.com', 'www.elfuturodelpasado.com', 'www.com', 'books.google.com', 'www.atkearney.com', 'tribune.com', 'www.gfkamerica.com', 'britannica.com', 'www.com', 'books.google.com', 'www.nytimes.com', 'www.mercurynews.com', 'ar-tour.com', 'auditorium.com', 'books.google.com', 'books.google.com', 'geography.about.com', 'edition.cnn.com', 'roundtheworldmagazin.com', 'demographia.com', 'www.arwu.org', 'esa.un.org', 'www.worldhistory.org', 'olympic.org', 'whc.unesco.org', 'www.archaeology.org', 'seatemperature.org', 'romaperkyoto.org', 'www.metmuseum.org', 'www.laphamsquarterly.org', 'catholic-hierarchy.org', 'www.arwu.org', 'newadvent.org', 'catalog.hathitrust.org', 'www.pbs.org', 'newadvent.org', 'romanculture.org', 'cwur.org', 'www.pnac.org', 'wayback.archive-it.org', 'www.npr.org', 'observatoribarcelona.org', 'www.npr.org', 'newadvent.org', 'www.port-of-rome.org', 'www.pbs.org', 'www.nationalgeographic.org', ['the classical review '], ['european journal of political theory '], ['the american journal of philology '], ['classical philology ', 'university of chicago press '], ['international journal of urban and regional research '], ['antiquity ', 'cambridge university press ']]",25458,Require autoconfirmed or confirmed access (no expiry set),203390,13 October 2001,BenBaker ,11705,18,2001-10-13,2001-10,2001
200,200,Greenland,https://en.wikipedia.org/wiki/Greenland,196,15,"['10.1086/303038', '10.1111/j.1751-8369.1997.tb00252.x', '10.1016/j.ajhg.2014.11.012', '10.3402/ijch.v71i0.18444', '10.1080/00438243.1999.9980423', '10.1029/96eo00142', '10.1093/biosci/bix014', '10.1080/03468750701449554', '10.3402/ijch.v72i0.19558', '10.3368/aa.50.1.72', '10.1525/aa.1940.42.3.02a00080', '10.1080/0108464x.1988.10589995', '10.1073/pnas.0902522107', '10.3721/037.002.s206', '10.3402/ijch.v64i3.17987', '10924403', None, '25557782', '23256091', None, None, '28608869', None, '23431117', None, None, None, '20212157', None, '16050317', '1287530', None, '4289681', '3525923', None, None, '5451287', None, '3577920', None, None, None, '2851789', None, None]","[['american journal of human genetics '], ['polar research '], ['american journal of human genetics '], ['international journal of circumpolar health '], ['world archaeology '], ['eos'], ['bioscience'], ['scandinavian journal of history ', 'scandinavian journal of history volume 33'], ['int j circumpolar health '], ['arctic anthropology '], ['american anthropologist '], ['journal of danish archaeology '], ['proceedings of the national academy of sciences '], ['journal of the north atlantic '], ['international journal of circumpolar health ']]",15,4,1,57,0,2,102,0.07653061224489796,0.02040816326530612,0.29081632653061223,0.07653061224489796,0.00510204081632653,0.17857142857142858,15,"['www.cia.gov', 'www.cia.gov', 'cia.gov', 'www.cia.gov', 'www.fodors.com', 'dotearth.blogs.nytimes.com', 'stalvik.com', 'books.google.com', 'www.airgreenland.com', 'ancientstandard.com', 'blogs.aljazeera.com', 'news.nationalgeographic.com', 'greenland.com', 'www.businessinsider.com', 'www.airgreenland.com', 'books.google.com', 'www.smithsonianmag.com', 'www.greenland.com', 'greenland.com', 'www.cbsnews.com', 'www.bbc.com', 'ams.confex.com', 'greenland.com', 'canada.com', 'books.google.com', 'greenland.com', 'news.nationalgeographic.com', 'www.nytimes.com', 'www.time.com', 'www.greenland.com', 'jazbablog.com', 'blog.oup.com', 'www.nytimes.com', 'www.theaustralian.news.com', 'www.businessweek.com', 'books.google.com', 'books.google.com', 'www.weather-atlas.com', 'www.washingtonpost.com', 'andrewskurth.com', 'thearda.com', 'www.arctictoday.com', 'news.google.com', 'www.greenland.com', 'books.google.com', 'books.google.com', 'www.wendyperrin.com', 'www.economist.com', 'news.nationalgeographic.com', 'www.nationaljeweler.com', 'books.google.com', 'www.iexplore.com', 'www.foxnews.com', 'www.smithsonianmag.com', 'www.cntraveler.com', 'worldislandinfo.com', 'www.nytimes.com', 'www.vice.com', 'books.google.com', 'www.slate.com', 'www.nationalreview.com', 'www.pewforum.org', 'www.operationworld.org', 'data.worldbank.org', 'data.worldbank.org', 'www.icj-cij.org', 'www.americanscientist.org', 'www.nautilus.org', 'www.nordiclabourjournal.org', 'data.worldbank.org', 'www.cidob.org', 'www.archaeology.org', 'unstats.un.org', 'www.thearcticinstitute.org', 'gutenberg.org', 'www.oikoumene.org', ['american journal of human genetics '], ['polar research '], ['american journal of human genetics '], ['international journal of circumpolar health '], ['world archaeology '], ['eos'], ['bioscience'], ['scandinavian journal of history ', 'scandinavian journal of history volume 33'], ['int j circumpolar health '], ['arctic anthropology '], ['american anthropologist '], ['journal of danish archaeology '], ['proceedings of the national academy of sciences '], ['journal of the north atlantic '], ['international journal of circumpolar health ']]",12118,Require administrator access (no expiry set),152102,4 May 2001,KoyaanisQatsi ,7355,2,2001-05-04,2001-05,2001
201,201,Eritrea,https://en.wikipedia.org/wiki/Eritrea,228,3,"['10.1126/science.1078208', '10.1038/35011048', '10.2307/1357309', '12714734', '10811218', None, None, None, None]","[[' science '], [' nature '], ['bulletin of the american schools of oriental research']]",52,4,0,101,0,8,60,0.22807017543859648,0.017543859649122806,0.44298245614035087,0.013157894736842105,0.0,0.25877192982456143,3,"['www.cia.gov', 'www.uscirf.gov', 'www.cia.gov', '2009-2017.state.gov', 'edition.cnn.com', 'dankalia.com', 'www.bloomberg.com', 'www.caperi.com', 'utdailybeacon.com', 'www.newsweek.com', 'www.procyclingstats.com', 'www.nytimes.com', 'books.google.com', 'books.google.com', 'www.addistribune.com', 'workmall.com', 'comstat.com', 'www.shabait.com', 'dictionary.com', 'www.washingtonpost.com', 'www.google.com', 'www.google.com', 'www.shabait.com', 'www.embassy-worldwide.com', 'www.google.com', 'thediplomat.com', 'books.google.com', 'www.voanews.com', 'www.weatherbase.com', 'books.google.com', 'books.google.com', 'allafrica.com', 'www.sudantribune.com', 'www.fatbirder.com', 'www.sudantribune.com', 'shabait.com', 'dadfeatured.blogspot.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'www.eritreanbeauty.com', 'books.google.com', 'shabait.com', 'www.washingtoncitypaper.com', 'dw.com', 'www.ethnologue.com', 'britannica.com', 'www.google.com', 'af.reuters.com', 'www.africanews.com', 'www.google.com', 'www.economist.com', 'www.addistribune.com', 'qz.com', 'shabait.com', 'eri24.com', 'www.aljazeera.com', 'books.google.com', 'www.bbc.com', 'www.voanews.com', 'www.freeourparents-eritrea.com', 'books.google.com', 'cqranking.com', 'www.google.com', 'www.statoids.com', 'www.madote.com', 'www.mining-technology.com', 'bloomberg.com', 'raimoq.com', 'smh.com', 'books.google.com', 'ibis.atwebpages.com', 'www.google.com', 'books.google.com', 'ibis.atwebpages.com', 'books.google.com', 'www.shabait.com', 'www.bbc.com', 'www.networkafricaonline.com', 'www.google.com', 'www.dw.com', 'www.sbs.com', 'www.google.com', 'www.caperi.com', 'books.google.com', 'books.google.com', 'washingtontimes.com', 'raimoq.com', 'www.google.com', 'www.nytimes.com', 'books.google.com', 'globaltwitcher.com', 'books.google.com', 'www.smithsonianmag.com', 'www.apollo-magazine.com', 'shabait.com', 'www.dw.com', 'www.voanews.com', 'books.google.com', 'www.washingtonpost.com', 'books.google.com', 'www.huffingtonpost.com', 'www.cyclingnews.com', 'explore-eritrea.com', 'www.google.com', 'www.imf.org', 'www.viv-it.org', 'daccess-dds-ny.un.org', 'www.fao.org', 'www.pewforum.org', 'www.pewresearch.org', 'whc.unesco.org', 'afdb.org', 'www.worldhistory.org', 'www.dskmariam.org', 'beta.thegef.org', 'en.rsf.org', 'rsf.org', 'www.iso.org', 'www.africabib.org', 'www.trainweb.org', 'population.un.org', 'www.irinnews.org', 'www.ohchr.org', 'databank.worldbank.org', 'www.odi.org', 'www.wri-irg.org', 'www.ohchr.org', 'www.hrw.org', 'uis.unesco.org', 'whc.unesco.org', 'uis.unesco.org', 'data.worldbank.org', 'www.unicef.org', 'dacb.org', 'www.nyulawglobal.org', 'er.undp.org', 'rsf.org', 'meeting.physanth.org', 'www.hrw.org', 'globalreligiousfutures.org', 'www.shaebia.org', 'www.hrw.org', 'hdr.undp.org', 'www.grassrootsonline.org', 'hrc-eritrea.org', 'imf.org', 'thebestofafrica.org', 'www.cpj.org', 'www.ehrea.org', 'jw.org', 'jw.org', 'www.worldbank.org', 'shaebia.org', 'www.africabib.org', 'www.unesco.org', 'iaaf.org', [' science '], [' nature '], ['bulletin of the american schools of oriental research']]",17238590,"Require autoconfirmed or confirmed access (16:47, 6 May 2023)",147826,30 September 2001,Ap ,8654,35,2001-09-30,2001-09,2001
202,202,Ukraine,https://en.wikipedia.org/wiki/Ukraine,454,15,"['10.3138/9781442682252', '10.18647/2730/jjs-2007', '10.1093/past/179.1.197', '10.1371/journal.pone.0020834', '10.1080/00085006.2007.11092432', '10.2307/3650068', '10.3390/su9071152', '10.1093/biosci/bix014', '10.1080/00905990500193204', '10.2307/1149308', '10.1111/1758-5899.12301', '10.1016/j.ejrh.2020.100761', '10.12911/22998993/132945', None, None, None, None, None, None, None, '28608869', None, None, None, None, None, None, None, None, None, None, None, None, '5451287', None, None, None, None, None]","[['university of toronto press '], ['the journal of jewish studies '], ['past '], ['plos one ', 'plos one '], ['canadian slavonic papers '], ['slavic review '], [' sustainability '], ['bioscience '], ['nationalities papers '], ['[[foreign policy'], ['[[global policy'], ['journal of hydrology'], ['journal of ecological engineering ']]",82,44,0,204,0,12,101,0.18061674008810572,0.09691629955947137,0.44933920704845814,0.03303964757709251,0.0,0.31057268722466963,13,"['www.mfa.gov', 'peremoga.gov', 'ukrcensus.gov', 'export.gov', 'www.state.gov', 'zakon1.rada.gov', 'www.education.gov', 'rv.gov', 'gska2.rada.gov', '2001.ukrcensus.gov', 'gska2.rada.gov', '2001-2009.state.gov', 'www.mil.gov', '2001.ukrcensus.gov', 'permanent.access.gpo.gov', 'peremoga.gov', 'www.archives.gov', 'portal.rada.gov', 'gska2.rada.gov', 'www.ukrstat.gov', 'www.cia.gov', 'peremoga.gov', 'moz.gov', 'ukrcensus.gov', 'www.cvk.gov', 'ukraineinvest.gov', 'www.mil.gov', 'gska2.rada.gov', 'www.nrada.gov', 'mvs.gov', 'www.education.gov', 'zakon.rada.gov', 'www.mil.gov', 'bank.gov', 'www.kmu.gov', 'www.derzhkomrelig.gov', 'www.mil.gov', 'zakon1.rada.gov', 'www.nkau.gov', 'ukrcensus.gov', '2009-2017.state.gov', 'w1.c1.rada.gov', 'www.cia.gov', 'education.gov', 'www.nytimes.com', 'www.nytimes.com', 'www.nytimes.com', 'www.bbc.com', 'en.interfax.com', 'www.nytimes.com', 'www.britannica.com', 'www.bbc.com', 'www.nytimes.com', 'www.wsj.com', 'www.kyivpost.com', 'birdinflight.com', 'ukrainianweek.com', 'www.euronews.com', 'www.kyivpost.com', 'books.google.com', 'life.pravda.com', 'for-ua.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'findarticles.com', 'www.bartleby.com', 'books.google.com', 'www.britannica.com', 'www.kyivpost.com', 'books.google.com', 'www.reuters.com', 'www.pravda.com', 'newlinesmag.com', 'books.google.com', 'www.britannica.com', 'www.themoscowtimes.com', 'books.google.com', 'www.routesonline.com', 'europe-cities.com', 'www.nytimes.com', 'www.ukraine.com', 'www.kyivpost.com', 'www.bloomberg.com', 'www.euractiv.com', 'www.britannica.com', 'www.usnews.com', 'kiis.com', 'archunion.com', 'www.mentalfloss.com', 'www.reuters.com', 'www.kyivpost.com', 'books.google.com', 'encyclopediaofukraine.com', 'www.washingtonpost.com', 'www.encyclopediaofukraine.com', 'www.pravda.com', 'www.dw.com', 'www.encyclopediaofukraine.com', 'www.ukrweekly.com', 'books.google.com', 'books.google.com', 'www.encyclopediaofukraine.com', 'www.reuters.com', 'nbnews.com', 'vicenews.com', 'books.google.com', 'www.vivafitness.com', 'apnews.com', 'books.google.com', 'www.britannica.com', 'slate.com', 'www.encyclopediaofukraine.com', 'www.nybooks.com', 'www.upi.com', 'www.newsweek.com', 'www.encyclopediaofukraine.com', 'ua-travelling.com', 'www.kyivpost.com', 'books.google.com', 'ukraine.com', 'www.ukrweekly.com', 'ndtv.com', 'encarta.msn.com', 'www.kyivpost.com', 'ukrferry.com', 'www.irishtimes.com', 'books.google.com', 'www.nybooks.com', 'books.google.com', 'www.foxnews.com', '(kiis.com', 'www.aljazeera.com', 'kyivpost.com', 'books.google.com', 'www.wsj.com', 'www.ukraine-observer.com', 'books.google.com', 'www.wsj.com', 'trackandfieldnews.com', 'www.reuters.com', 'www.reuters.com', 'www.reuters.com', 'www.aljazeera.com', 'religiya_200516_a4.com', 'www.economist.com', 'www.britannica.com', 'www.usatoday.com', 'www.cbsnews.com', 'en.for-ua.com', 'books.google.com', 'www.nytimes.com', 'www.thedailybeast.com', 'www.wsj.com', 'www.britannica.com', 'www.sciencedaily.com', 'www.businessinsider.com', 'www.bbc.com', 'www.nytimes.com', 'www.britannica.com', 'www.britannica.com', 'www.bloombergquint.com', 'www.cbsnews.com', 'www.schengenvisainfo.com', 'www.nytimes.com', 'www.britannica.com', 'www.nytimes.com', 'www.kyivpost.com', 'www.britannica.com', 'www.ceicdata.com', 'www.whichairline.com', 'www.kyivpost.com', 'www.nytimes.com', 'www.pravda.com', 'books.google.com', 'kyivpost.com', 'www.flyuia.com', 'www.kyivpost.com', 'europeanvoice.com', 'www.nytimes.com', 'religiya_200516_a4.com', '(www.dw.com', 'apnews.com', 'ndtv.com', 'kyivpost.com', 'www.rlef.eu.com', 'www.tourismroi.com', 'www.merriam-webster.com', 'books.google.com', 'www.theatlantic.com', 'businessweek.com', 'www.nytimes.com', 'www.nytimes.com', 'www.kyivpost.com', 'nytimes.com', 'www.eurointegration.com', 'radiolemberg.com', 'www.nytimes.com', 'dw.com', 'theconversation.com', 'www.britannica.com', 'www.euractiv.com', 'books.google.com', 'uk.reuters.com', 'www.britannica.com', 'www.westinghousenuclear.com', 'www.dailykos.com', 'cbsnews.com', 'cnn.com', 'books.google.com', 'apnews.com', 'encyclopediaofukraine.com', 'en.interfax.com', 'en.interfax.com', 'emerging-europe.com', 'en.interfax.com', 'www.nytimes.com', 'www.britannica.com', 'www.economist.com', 'www.nytimes.com', 'books.google.com', 'www.businessukraine.com', 'www.bbc.com', 'britannica.com', 'books.google.com', 'www.encyclopediaofukraine.com', 'ukranews.com', 'rb.com', 'www.ft.com', 'www.bbc.com', 'www.encyclopediaofukraine.com', 'topics.nytimes.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'www.ft.com', 'www.ditext.com', 'books.google.com', 'www.bbc.com', 'www.economist.com', 'bbcukrainian.com', 'www.kyivpost.com', 'www.euronews.com', 'bestofukraine.com', 'global.britannica.com', 'www.britannica.com', 'espn.com', 'www.worldbank.org', 'data.worldbank.org', 'climateknowledgeportal.worldbank.org', 'ukrstat.org', 'www.atlanticcouncil.org', 'niisp.org', 'razumkov.org', 'data.worldbank.org', 'imf.org', 'www.transparency.org', 'www.jstor.org', 'freedomhouse.org', 'www.imf.org', 'usva.org', 'www.ramsar.org', 'imf.org', 'www.ramsar.org', 'www.un.org', 'data2.unhcr.org', 'www.jamestown.org', 'www.worldbank.org', 'www.fao.org', 'www.worldcat.org', 'norric.org', 'unesdoc.unesco.org', 'ti-ukraine.org', 'www.hrw.org', 'www.migrationpolicy.org', 'www.rferl.org', 'www.pewforum.org', 'ceobs.org', 'translatorswithoutborders.org', 'whc.unesco.org', 'www.radiosvoboda.org', 'preferredbynature.org', 'www.rferl.org', 'voxukraine.org', 'www.imf.org', 'www.unicef.org', 'old.razumkov.org', 'ich.unesco.org', 'www.osce.org', 'en.wikisource.org', 'www.oecd-ilibrary.org', 'whc.unesco.org', 'www.atlanticcouncil.org', 'uacrisis.org', 'data.worldjusticeproject.org', 'www.un.org', 'www.jamestown.org', 'old.razumkov.org', 'data.worldbank.org', 'www.pewforum.org', 'www.nti.org', 'www.jstor.org', 'www.unicef.org', 'www.fao.org', 'warhistory.ukrlife.org', 'www.rferl.org', 'freedomhouse.org', 'ich.unesco.org', 'www.osce.org', 'fas.org', 'devdata.worldbank.org', 'uacrisis.org', 'openknowledge.worldbank.org', 'imh.org', 'www.olympic.org', 'www.fao.org', 'ich.unesco.org', 'www.npr.org', 'jamestown.org', 'www.iea.org', 'www.radiosvoboda.org', 'www.umacleveland.org', 'fmm51.org', 'hdr.undp.org', 'ukrstat.org', 'www.wto.org', 'www.iaea.org', 'www.iccrimea.org', 'globalsecurity.org', ['university of toronto press '], ['the journal of jewish studies '], ['past '], ['plos one ', 'plos one '], ['canadian slavonic papers '], ['slavic review '], [' sustainability '], ['bioscience '], ['nationalities papers '], ['[[foreign policy'], ['[[global policy'], ['journal of hydrology'], ['journal of ecological engineering ']]",31750,Require administrator access (no expiry set),263582,25 September 2001,195.206.85.xxx ,14143,99,2001-09-25,2001-09,2001
203,203,Cornwall,https://en.wikipedia.org/wiki/Cornwall,207,3,"['10.1017/s0079497x00000293', '10.1111/1469-8219.00027', '10.1371/journal.pone.0218326', None, None, '31242218', None, None, '6594607']","[[' proceedings of the prehistoric society', ' the prehistoric society'], [' nations and nationalism'], [' plos one ']]",25,22,0,39,0,1,117,0.12077294685990338,0.10628019323671498,0.18840579710144928,0.014492753623188406,0.0,0.24154589371980675,3,"['www.gov', 'www.cornwall.gov', 'www.cornwall.gov', 'www.cornwall.gov', 'www.scottishexecutive.gov', 'www.gov', 'www.metoffice.gov', 'www.cornwall-aonb.gov', 'www.cornwall.gov', 'www.cornwall.gov', 'db.cornwall.gov', 'www.onecornwall.cornwall.gov', 'wales.gov', 'www.cornwall.gov', 'www.gov', 'www.cornwall.gov', 'www.cornwall.gov', 'www.ons.gov', 'www.ons.gov', 'www.ons.gov', 'www.cornwall.gov', 'www.cornwall.gov', 'books.google.com', 'oxforddictionaries.com', 'www.visitcornwall.com', 'www.oxbowbooks.com', 'www.channel4.com', 'crwflags.com', 'www.etymonline.com', 'www.metoffice.com', 'southwestcoastpath.com', 'thefreedictionary.com', 'www.etymonline.com', 'www.nytimes.com', 'books.google.com', 'www.moviediva.com', 'third-millennium-library.com', 'books.google.com', 'glosbe.com', 'www.theage.com', 'www.cprw.com', 'www.visitcornwall.com', 'www.artnet.com', 'severnlink.com', 'www.metoffice.com', 'www.festival-interceltique.com', 'www.authorama.com', 'submarinecablemap.com', 'www.stormfinearts.com', 'www.st-piran.com', 'datasegment.com', 'www.oxforddnb.com', 'www.marketwired.com', 'www.metoffice.com', 'www.cornwalllive.com', 'an-daras.com', 'www.powells.com', 'www.studio-pots.com', 'dailyhomelist.com', 'edition.cnn.com', 'objectiveone.com', 'welshjournals.llgc.org', 'visionofbritain.org', 'www.flaginstitute.org', 'visionofbritain.org', 'www.superfastcornwall.org', 'www.penleehouse.org', 'www.hp-lexicon.org', 'www.worldwideschool.org', 's-gabriel.org', 'www.celtic-congress.org', 'www.dumaurier.org', 'whc.unesco.org', 'linecaught.org', 'www.tate.org', 'www.plymouth-diocese.org', 'www.trurocathedral.org', '.org', 'www.mebyonkernow.org', 'cornwallstatistics.org', 'cornish-mining.org', 'alanrichards.org', 'cornishassembly.org', 'www.cornish-mining.org', 'newlynfishfestival.org', 'cornishassembly.org', [' proceedings of the prehistoric society', ' the prehistoric society'], [' nations and nationalism'], [' plos one ']]",5648,Allow all users (no expiry set),140986,12 October 2001,J Hofmann Kemp ,6404,17,2001-10-12,2001-10,2001
204,204,Hyderabad,https://en.wikipedia.org/wiki/Hyderabad,355,6,"['10.1080/13602008508715945', '10.1017/s0026749x00004996', '10.1080/19472498.2011.577568', '10.3390/ijerph2005020021', '10.1136/ip.2008.019620', '10.1080/02666030.1993.9628458', None, None, None, '16705838', '19074239', None, None, None, None, '3810641', '2777413', None]","[['journal of muslim minority affairs '], ['[[modern asian studies'], ['south asian history and culture '], ['international journal of environmental research and public health '], ['injury prevention '], ['south asian studies ']]",27,38,0,186,0,0,98,0.07605633802816901,0.10704225352112676,0.523943661971831,0.016901408450704224,0.0,0.2,6,"['www.mhrd.gov', 'www.hyderabadwater.gov', 'ccrtindia.gov', 'www.ded.mo.gov', 'ghmc.gov', 'www.aponline.gov', 'hyderabadpolice.gov', 'www.ghmc.gov', 'cgg.gov', 'scb.aponline.gov', 'aponline.gov', 'www.apdes.ap.gov', 'www.imdhyderabad.gov', 'aponline.gov', 'pdf.usaid.gov', 'www.cyberabadpolice.gov', 'aponline.gov', 'www.apind.gov', 'www.censusindia.gov', 'www.delhi.gov', 'pdf.usaid.gov', 'www.ghmc.gov', 'censusindia.gov', 'www.scr.indianrailways.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'aponline.gov', 'aponline.gov', 'www.imd.gov', 'cgg.gov', 'www.censusindia.gov', 'www.hmda.gov', 'invest.telangana.gov', 'www.forests.ap.gov', 'www.cia.gov', 'www.ghmc.gov', 'www.ghmc.gov', 'www.ghmc.gov', 'www.ndtv.com', 'rediff.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'hindu.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'www.hydzoo.com', 'www.thehindu.com', 'www.thehindu.com', 'www.hindu.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.hindu.com', 'world.time.com', 'epaper.thehansindia.com', 'timesofindia.indiatimes.com', 'www.deccanchronicle.com', 'www.nytimes.com', 'www.news18.com', 'www.hindu.com', 'timesofindia.indiatimes.com', 'www.ndtv.com', 'www.deccanchronicle.com', 'www.newindianexpress.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.hindu.com', 'www.hindu.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'telanganatoday.com', 'timesofindia.indiatimes.com', 'articles.timesofindia.indiatimes.com', 'articles.timesofindia.indiatimes.com', 'www.livemint.com', 'timesofindia.indiatimes.com', 'www.livemint.com', 'www.deccanchronicle.com', 'books.google.com', 'www.thehindu.com', 'www.northbridgeasia.com', 'timesofindia.indiatimes.com', 'rediff.com', 'www.hyderabadliteraryfestival.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.greaterkashmir.com', 'www.thehindu.com', 'www.hindustantimes.com', 'books.google.com', 'ontheshortwaves.com', 'www.nytimes.com', 'timesofindia.indiatimes.com', 'ibnlive.in.com', 'www.business-standard.com', 'maps.google.com', 'www.livemint.com', 'timesofindia.indiatimes.com', 'www.milligazette.com', 'www.hindu.com', 'www.hindu.com', 'www.siasat.com', 'archives.deccanchronicle.com', 'www.thehindu.com', 'books.google.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'ibnlive.in.com', 'books.google.com', 'hindu.com', 'www.dnaindia.com', 'rediff.com', 'www.livemint.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'www.saudiaramcoworld.com', 'www.livemint.com', 'www.thehindu.com', 'www.publishersglobal.com', 'www.guinnessworldrecords.com', 'rediff.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'archive.indianexpress.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'rediff.com', 'www.thehindubusinessline.com', 'www.newindianexpress.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.hindu.com', 'timesofindia.indiatimes.com', 'archive.indianexpress.com', 'www.siasat.com', 'timesofindia.indiatimes.com', 'www.hindu.com', 'www.thehindu.com', 'www.tssouthernpower.com', 'www.thehindu.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.thehindu.com', 'postnoon.com', 'timesofindia.indiatimes.com', 'www.livemint.com', 'timesofindia.indiatimes.com', 'www.ukmediacentre.pwc.com', 'books.google.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'books.google.com', 'ibnlive.in.com', 'www.thehindu.com', 'www.siasat.com', 'www.thehindu.com', 'www.thehindu.com', 'www.livemint.com', 'timesofindia.indiatimes.com', 'jntuhdufr.com', 'www.deccanchronicle.com', 'www.hindu.com', 'www.hindu.com', 'timesofindia.indiatimes.com', 'www.huffingtonpost.com', 'timesofindia.indiatimes.com', 'www.siasat.com', 'timesofindia.indiatimes.com', 'www.hindu.com', 'www.thehindubusinessline.com', 'www.hindu.com', 'www.worldstadiums.com', 'www.hindu.com', 'www.hindu.com', 'www.hindu.com', 'books.google.com', 'books.google.com', 'careers.microsoft.com', 'www.docstoc.com', 'www.hindu.com', 'www.firstpost.com', 'www.worldstadiums.com', 'archive.indianexpress.com', 'hindu.com', 'www.weatherbase.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'www.weatherbase.com', 'timesofindia.indiatimes.com', 'books.google.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'indianexpress.com', 'timesofindia.indiatimes.com', 'www.hindu.com', 'insideismailism.files.wordpress.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehindu.com', 'www.hindu.com', 'www.livemint.com', 'www.deccanchronicle.com', 'www.thehindu.com', 'books.google.com', 'www.hindu.com', 'books.google.com', 'hindu.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.britishmuseum.org', 'siteresources.worldbank.org', 'www.itdp.org', 'www.unesco.org', 'saciwaters.org', 'www.unescobkk.org', 'jhss.org', 'en.unesco.org', 'prsindia.org', 'www.tnsroindia.org', 'www.redress.org', 'www.safewaternetwork.org', 'rainwaterharvesting.org', 'www.itdp.org', 'www.mciindia.org', 'circed.org', 'www.albioncx19project.org', 'www.un.org', 'cseindia.org', 'nasvinet.org', 'www.apeamcet.org', 'jointactionforwater.org', 'whc.unesco.org', 'indianheartassociation.org', 'www.doingbusiness.org', 'www.cicred.org', 'www.sundarayya.org', ['journal of muslim minority affairs '], ['[[modern asian studies'], ['south asian history and culture '], ['international journal of environmental research and public health '], ['injury prevention '], ['south asian studies ']]",37534,Require autoconfirmed or confirmed access (no expiry set),220021,3 February 2002,130.94.122.xxx ,16816,48,2002-02-03,2002-02,2002
205,205,Vikings,https://en.wikipedia.org/wiki/Vikings,326,17,"['10.1002/wea.150', '10.1227/01.neu.0000144825.92264.c4', '10.1093/molbev/msm255', '10.1002/9780470995501.ch7', '10.1002/ajpa.23308', '10.1016/j.evolhumbehav.2016.10.013', '10.1016/j.ehb.2019.05.007', '10.1034/j.1600-0390.2000.d01-1.x', '10.1016/j.jasrep.2017.02.014', '10.1111/j.1478-0542.2011.00820.x', '10.1002/ana.410360810', '10.1038/s41586-020-2688-8', '10.2307/2864557', '10.1179/007660905x54080', '10.1086/318785', '10.1484/j.jml.3.26', None, '16331154', '18032405', None, '28884802', None, '31208936', None, None, None, '7998792', '32939067', None, None, '11179019', None, None, None, '2628767', None, '5724682', None, None, None, None, None, None, None, None, None, '1274484', None]","[['weather'], ['neurosurgery '], ['molecular biology and evolution '], ['blackwell '], ['american journal of physical anthropology'], ['evolution and human behavior'], ['economics and human biology'], ['acta archaeologica'], ['journal of archaeological science'], ['history compass'], ['annals of neurology'], ['nature'], ['speculum'], ['medieval archaeology '], [' the american journal of human genetics'], ['the journal of medieval latin']]",18,3,0,96,0,1,191,0.05521472392638037,0.009202453987730062,0.294478527607362,0.05214723926380368,0.0,0.1165644171779141,16,"['lepel.vitebsk-region.gov', 'www.royal.gov', 'www.royal.gov', 'www.britannica.com', 'freya.theladyofthelabyrinth.com', 'www.livescience.com', 'books.google.com', 'blog.oup.com', 'www.britannica.com', 'www.forbes.com', 'www.nationalgeographic.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.straightdope.com', 'www.britannica.com', 'brill.com', 'books.google.com', 'archeurope.com', 'www.oed.com', 'books.google.com', 'www.oxbowbooks.com', 'www.wired.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.vikinganswerlady.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.cnn.com', 'books.google.com', 'www.historyextra.com', 'news.scotsman.com', 'www.etymonline.com', 'www.collinsdictionary.com', 'bunews.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.familytreedna.com', 'blogs.discovermagazine.com', 'www.livescience.com', 'www.smithsonianmag.com', 'www.youtube.com', 'books.google.com', 'books.google.com', 'muslimheritage.com', 'www.destructoid.com', 'www.livescience.com', 'archive.aramcoworld.com', 'news.nationalgeographic.com', 'www.economist.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'dictionary.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'www.nature.com', 'brill.com', 'books.google.com', 'www.gameinformer.com', 'www.thevintagenews.com', 'books.google.com', 'books.google.com', 'books.google.com', 'sciencenordic.com', 'books.google.com', 'www.oxfordreference.com', 'www.oxfordreference.com', 'www.scribd.com', 'books.google.com', 'realscandinavia.com', 'www.collinsdictionary.com', 'books.google.com', 'vasmer.slovaronline.com', 'www.smithsonianmag.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.encyclopediaofukraine.com', 'books.google.com', 'www.nbcnews.com', 'books.google.com', 'books.google.com', 'sciencenordic.com', 'www.sciencealert.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.britannica.com', 'docs.wixstatic.com', 'www.collinsdictionary.com', 'dougcabot.com', 'allthatsinteresting.com', 'books.google.com', 'archive.archaeology.org', 'dictionary.cambridge.org', 'www.sciencemag.org', 'metmuseum.org', 'www.sciencemag.org', 'www.archaeology.org', 'www.archaeology.org', 'www.hoover.org', 'www.sciencemag.org', 'dragonslaire.org', 'www.sciencemag.org', 'www.pbs.org', 'nvg.org', 'www.regia.org', 'www.sciencemag.org', 'runeberg.org', 'runeberg.org', 'www.worldhistory.org', ['weather'], ['neurosurgery '], ['molecular biology and evolution '], ['blackwell '], ['american journal of physical anthropology'], ['evolution and human behavior'], ['economics and human biology'], ['acta archaeologica'], ['journal of archaeological science'], ['history compass'], ['annals of neurology'], ['nature'], ['speculum'], ['medieval archaeology '], [' the american journal of human genetics'], ['the journal of medieval latin']]",32610,Require autoconfirmed or confirmed access (no expiry set),196629,16 October 2001,Sjc ,7646,2,2001-10-16,2001-10,2001
206,206,Spain,https://en.wikipedia.org/wiki/Spain,320,9,"['10.1126/science.1219957', '10.1136/bmj.n1343', '10.1163/9789004443594_006', '10.1177/23409444211042382', '10.26882/histagrar.083e08p', '10.15304/9788416533015', '10.1038/s41467-020-19493-3', '10.1093/reseval/rvaa014', '10.1515/9783110365955-018', '22700921', '34162598', None, None, None, None, '33293507', None, None, None, '8220857', None, None, None, None, '7723057', None, None]","[['science'], ['bmj'], ['[[brill '], ['business research quarterly'], ['historia agraria'], ['servizo de publicacións e intercambio científico da universidade de compostela'], ['nature communications'], ['research evaluation'], ['[[de gruyter']]",42,8,0,104,0,6,152,0.13125,0.025,0.325,0.028125,0.0,0.184375,9,"['www.fco.gov', 'lcweb2.loc.gov', 'lcweb2.loc.gov', 'www.cia.gov', 'lcweb2.loc.gov', 'lcweb2.loc.gov', 'lcweb2.loc.gov', 'cia.gov', 'www.iht.com', 'books.google.com', 'www.economist.com', 'books.google.com', 'www.trobat.com', 'elpais.com', 'books.google.com', 'blogs.wsj.com', 'www.bbc.com', 'books.google.com', 'www.elperiodico.com', 'worldpridemadrid2017.com', 'justiciadegenero.com', 'www.economist.com', 'www.elpais.com', 'www.lavanguardia.com', 'noticias.juridicas.com', 'leekuanyewworldcityprize.com', 'elpais.com', 'bloomberg.com', 'www.elespanol.com', 'www.newscientist.com', 'www.economist.com', 'thehistorynet.com', 'www.washingtonpost.com', 'www.economist.com', 'www.economist.com', 'books.google.com', 'workpermit.com', 'www.bbc.com', 'www.economist.com', 'www.wsj.com', 'books.google.com', 'www.audiovisual451.com', 'www.elpais.com', 'www.economist.com', 'www.businessweek.com', 'www.economist.com', 'books.google.com', 'elpais.com', 'politica.elpais.com', 'www.iht.com', 'www.wsj.com', 'www.theglobalguru.com', 'linguatics.com', 'www.economist.com', 'books.google.com', 'books.google.com', 'books.google.com', 'elpais.com', 'books.google.com', 'books.google.com', 'europeanfutureenergyforum.com', 'www.forbes.com', 'elpais.com', 'www.demographia.com', 'books.google.com', 'noticias.juridicas.com', 'www.statista.com', 'triplepundit.com', 'www.theportugalnews.com', 'elpais.com', 'city-data.com', 'www.nytimes.com', 'books.google.com', 'www.moroccoworldnews.com', 'books.google.com', 'books.google.com', 'www.euronews.com', 'triplepundit.com', 'encarta.msn.com', 'worldmayor.com', 'books.google.com', 'learnodo-newtonic.com', 'www.theglobalguru.com', 'www.scimagoir.com', 'www.elpais.com', 'noticias.juridicas.com', 'books.google.com', 'edition.cnn.com', 'books.google.com', 'www.villagevoice.com', 'elpais.com', 'www.reuters.com', 'www.britannica.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'www.lavanguardia.com', 'blog.raileurope.com', 'books.google.com', 'bank-holidays.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'justiciadegenero.com', 'books.google.com', 'www.bbc.com', 'es.euronews.com', 'www.economist.com', 'www.channel4.com', 'www.theatlantic.com', 'www.msnbc.msn.com', 'ferede.org', 'upload.wikimedia.org', 'esa.un.org', 'www.un.org', 'data.worldbank.org', 'stats.oecd.org', 'whc.unesco.org', 'www1.worldbank.org', 'www.unesco.org', 'www.redalyc.org', 'www.oecd.org', 'www.oecd.org', 'ourworldindata.org', 'churchofjesuschrist.org', 'imf.org', 'www2.compareyourcountry.org', 'www.osce.org', 'npr.org', 'www.worldvaluessurvey.org', 'daccess-dds-ny.un.org', 'hdr.undp.org', 'www1.worldbank.org', 'daccess-dds-ny.un.org', 'phys.org', 'www.eolicenergynews.org', 'ipu.org', 'www.oecd.org', 'www.jewishvirtuallibrary.org', 'www.aeeolica.org', 'www.earthtimes.org', 'hdr.undp.org', 'www.amnesty.org', 'www.un.org', 'cartujo.org', 'www.investinspain.org', 'www.pewglobal.org', 'www.eumap.org', 'www.movimientoeuropeo.org', 'www.understandinganimalresearch.org', '.gobiernodecanarias.org', 'www.eumap.org', 'www.cyberistan.org', ['science'], ['bmj'], ['[[brill '], ['business research quarterly'], ['historia agraria'], ['servizo de publicacións e intercambio científico da universidade de compostela'], ['nature communications'], ['research evaluation'], ['[[de gruyter']]",26667,Require administrator access (no expiry set),254432,3 October 2001,Tezcatlipoca ,16042,38,2001-10-03,2001-10,2001
207,207,Netherlands,https://en.wikipedia.org/wiki/Netherlands,311,8,"['10.1038/s41467-020-19493-3', '10.1177/0021140019872340', '10.1086/650185', '10.1073/pnas.1112261109', '10.1111/1539-6924.00338', '10.3390/resources7030058', '10.1038/466170a', '10.1093/biosci/bix014', '33293507', None, None, '22308348', '12836850', None, '20613812', '28608869', '7723057', None, None, '3277516', None, None, None, '5451287']","[['nature communications'], [' irish theological quarterly'], ['crime and justice'], ['proceedings of the national academy of sciences'], ['risk analysis '], ['resources'], ['nature'], ['bioscience']]",32,13,0,81,0,1,176,0.10289389067524116,0.04180064308681672,0.2604501607717042,0.02572347266881029,0.0,0.17041800643086816,8,"['www.cia.gov', 'www.fas.usda.gov', 'www.gov', 'cia.gov', 'cia.gov', 'www.gov', 'cia.gov', 'www.gov', 'factfinder.census.gov', 'lcweb2.loc.gov', 'www.cia.gov', '2009-2017.state.gov', 'www.cia.gov', 'worldatlas.com', 'books.google.com', 'books.google.com', 'healthpowerhouse.com', 'books.google.com', 'www.dutchdailynews.com', 'books.google.com', 'www.canto-ostinato.com', 'www.britannica.com', 's3.amazonaws.com', 'www.britannica.com', 'www.portofrotterdam.com', 'www.theverge.com', 'books.google.com', 'www.reuters.com', 'www.bbc.com', 'www.geoexpro.com', 'link.galegroup.com', 'books.google.com', 'www.netherlands-tourism.com', 'books.google.com', 'www.economist.com', 'books.google.com', 'www.forbes.com', 'hollandtrade.com', 'www.nytimes.com', 'www.nationalgeographic.com', 'www.boston.com', 'www.reuters.com', 'books.google.com', 'www.annualreportschiphol.com', 'necrometrics.com', 'local-life.com', 'books.google.com', 'books.google.com', 'happiness-report.s3.amazonaws.com', 'www.ibtimes.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'www.boston.com', 'www.france24.com', 'marketwatch.com', 'transcripts.cnn.com', 'allmusic.com', 'www.holland.com', 'about.com', 'www.ecf.com', 'www.encyclopedia.com', 'www.nwaonline.com', 'books.google.com', 'archiver.rootsweb.ancestry.com', 'hollandtrade.com', 'healthpowerhouse.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.forbes.com', 'dannyreviews.com', 'topics.nytimes.com', 'sustainablecitiesindex.com', 'www.billboard.com', 'channelnewsasia.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'edition.cnn.com', 'press.andrerieu.com', 'www.ft.com', 'books.google.com', 'www.consoglobe.com', 'www.bbc.com', 'books.google.com', 'www.allmusic.com', 'uk.reuters.com', 'handbook.reuters.com', 'www.freshplaza.com', 'www.britannica.com', 'www.timeanddate.com', 'www2.deloitte.com', 'www.news18.com', 'ourworldindata.org', 'www.iea.org', 'www.oxfamamerica.org', 'livius.org', 'de.scientificcommons.org', 'www.imd.org', 'npr.org', 'www.iea.org', 'repositories.cdlib.org', 'unicef-irc.org', 'www.ibiblio.org', 'www.imf.org', 'www.iea.org', 'news.sciencemag.org', 'internationaltransportforum.org', 'asce.org', 'www.iea.org', 'www.iea.org', 'nl.wikisource.org', 'netherlandsmission.org', 'www.heritage.org', 'content.healthaffairs.org', 'www.livius.org', 'beleven.org', 'rsf.org', 'data.footprintnetwork.org', 'data.worldbank.org', 'unicef.org', 'www.weforum.org', 'heritage.org', 'www.imf.org', 'hdr.undp.org', ['nature communications'], [' irish theological quarterly'], ['crime and justice'], ['proceedings of the national academy of sciences'], ['risk analysis '], ['resources'], ['nature'], ['bioscience']]",21148,Require administrator access (no expiry set),269989,15 November 2001,Stephen Gilbert ,17050,7,2001-11-15,2001-11,2001
208,208,Luo people,https://en.wikipedia.org/wiki/Luo_people,81,23,"['10.1371/journal.pgen.1006976', '10.1017/s0021853700021289', '10.1007/bf02860055', '10.2307/3556798', '10.1017/s002185370002973x', '10.1163/19589514-047-01-900000010', '10.2307/217849', '10.2307/3052969', '10.1126/science.1172257', '10.1080/00672700609480438', '10.2307/1581402', '10.1017/s0021853700010859', '10.2307/3097285', '10.1017/s0021853700027572', '10.1080/00672700903291716', '10.1086/201823', '10.1023/a:1019954903395', '10.21504/amj.v5i3.1658', '10.5070/d64110028', '10.1038/sj.ejhg.5201408', '10.1525/nr.2009.13.1.11', '10.1080/01436590120084575', '28837655', None, None, None, None, None, None, None, '19407144', None, None, None, None, None, None, None, None, None, None, '15856073', None, None, '5587336', None, None, None, None, None, None, None, '2947357', None, None, None, None, None, None, None, None, None, None, None, None, None]","[['plos genetics '], ['the journal of african history '], ['economic botany '], ['africa'], ['the journal of african history '], ['faits de langues '], ['the international journal of african historical studies '], ['law '], ['science '], ['azania'], ['journal of religion in africa '], ['the journal of african history '], ['the international journal of african historical studies '], ['the journal of african history '], ['azania'], ['current anthropology '], ['journal of world prehistory '], ['african music'], ['dotawo'], [' european journal of human genetics '], ['nova religio '], ['third world quarterly ']]",7,1,1,7,0,2,40,0.08641975308641975,0.012345679012345678,0.08641975308641975,0.2839506172839506,0.012345679012345678,0.3950617283950617,22,"['www.cia.gov', 'www.theafricareport.com', 'www.bbc.com', 'www.britannica.com', 'www.ethnologue.com', 'www.voanews.com', 'news.theage.com', 'www.newspapers.com', 'cotu-kenya.org', 'www.polity.org', 'www.amnesty.org', 'www.worldbank.org', 'nai.diva-portal.org', 'africanrockart.org', 'nai.diva-portal.org', ['plos genetics '], ['the journal of african history '], ['economic botany '], ['africa'], ['the journal of african history '], ['faits de langues '], ['the international journal of african historical studies '], ['law '], ['science '], ['azania'], ['journal of religion in africa '], ['the journal of african history '], ['the international journal of african historical studies '], ['the journal of african history '], ['azania'], ['current anthropology '], ['journal of world prehistory '], ['african music'], ['dotawo'], [' european journal of human genetics '], ['nova religio '], ['third world quarterly ']]",2771856,Allow all users (no expiry set),81347,26 September 2005,Ezeu ,1444,5,2005-09-26,2005-09,2005
209,209,Ladakh,https://en.wikipedia.org/wiki/Ladakh,146,6,"['10.1007/s00267-005-0178-2', '10.1111/j.1756-1051.2010.00983.x', '10.1007/s11284-006-0015-y', '10.1017/s0030605308000768', '10.1016/j.biocon.2005.09.003', '10.1007/s00267-005-0356-2', '17318699', None, None, None, None, '16955231', None, None, None, None, None, '1705511']","[['environmental management '], ['nordic journal of botany '], ['ecological research '], ['oryx '], ['biological conservation '], ['environmental management ']]",10,6,0,75,0,0,50,0.0684931506849315,0.0410958904109589,0.5136986301369864,0.0410958904109589,0.0,0.1506849315068493,6,"['results.eci.gov', 'allindiaradio.gov', 'www.ddindia.gov', 'www.censusindia.gov', 'censusindia.gov', 'dse.ladakh.gov', 'www.tribuneindia.com', 'books.google.com', 'www.britannica.com', 'timesofindia.indiatimes.com', 'www.jammu-kashmir.com', 'www.himalmag.com', 'www.oed.com', 'www.leh-ladakh-taxi-booking.com', 'books.google.com', 'ndtv.com', 'www.outlookindia.com', 'indianexpress.com', 'books.google.com', 'www.leh-ladakh-taxi-booking.com', 'www.thelalit.com', 'business-standard.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.dailyexcelsior.com', 'www.dollsofindia.com', 'www.powells.com', 'reachladakh.com', 'books.google.com', 'indianexpress.com', 'timesofindia.indiatimes.com', 'books.google.com', 'news.outlookindia.com', 'www.ndtv.com', 'www.greaterkashmir.com', 'books.google.com', 'peakbagger.com', 'www.nytimes.com', 'reference.allrefer.com', 'books.google.com', 'www.scmp.com', 'timesofindia.indiatimes.com', 'economictimes.indiatimes.com', 'books.google.com', 'www.business-standard.com', 'books.google.com', 'www.hindustantimes.com', 'books.google.com', 'ndtv.com', 'www.birdinginladakh.com', 'www.educationforallinindia.com', 'www.dailyexcelsior.com', 'www.scmp.com', 'books.google.com', 'www.amarujala.com', 'www.firstpost.com', 'lehladakhindia.com', 'www.dailyexcelsior.com', 'indianexpress.com', 'internationaledventures.com', 'www.thehindu.com', 'books.google.com', 'www.efi-news.com', 'www.economist.com', 'thaindian.com', 'indianexpress.com', 'books.google.com', 'www.thehindu.com', 'www.kashmirtimes.com', 'books.google.com', 'www.greaterkashmir.com', 'books.google.com', 'books.google.com', 'www.outlookindia.com', 'khagta.photoshelter.com', 'indianexpress.com', 'www.britannica.com', 'timesofindia.indiatimes.com', 'www.educationforallinindia.com', 'blog.cpsindia.org', 'www.jktourism.org', 'unesdoc.unesco.org', 'plantlife.org', 'www.hockeyfoundation.org', 'globalsecurity.org', 'wayback.archive-it.org', 'www.prsindia.org', 'www.icpsnet.org', 'www.universityofladakh.org', ['environmental management '], ['nordic journal of botany '], ['ecological research '], ['oryx '], ['biological conservation '], ['environmental management ']]",303611,Require autoconfirmed or confirmed access (no expiry set),115874,24 August 2003,Wik ,4060,9,2003-08-24,2003-08,2003
210,210,Traditional food,https://en.wikipedia.org/wiki/Traditional_food,40,3,"['10.14430/arctic1539', None, '10.1016/j.appet.2008.11.008', None, '7343324', '19084040', None, None, None]","[[' arctic'], ['food and agriculture organization of the united nations '], ['[[appetite ']]",1,0,0,28,0,0,8,0.025,0.0,0.7,0.075,0.0,0.1,3,"['visitcyprus.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'agriculturesociety.com', 'www.youtube.com', 'books.google.com', 'books.google.com', 'thezenchilada.com', 'books.google.com', 'www.bradenton.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.oxfordreference.com', 'www.afm-marketing.org', [' arctic'], ['food and agriculture organization of the united nations '], ['[[appetite ']]",46355870,Allow all users (no expiry set),31448,8 April 2015,Northamerica1000 ,412,0,2015-04-08,2015-04,2015
211,211,Iraq,https://en.wikipedia.org/wiki/Iraq,341,12,"['10.1093/biosci/bix014', '10.1007/s11159-005-0587-8', '10.1080/02684521003588120', '10.1163/157338410x12743419189540', '10.1038/srep04250', '10.1136/bmjgh-2017-000311', '10.1186/1471-2148-11-288', '10.1093/acref/9780195176322.001.0001', '10.2307/141771', '10.1515/libri-2015-0110', '28608869', None, None, None, '24603901', '29225933', '21970613', None, None, None, '5451287', None, None, None, '3945051', '5717930', '3215667', None, None, None]","[['bioscience'], ['international review of education'], ['intelligence and national security'], ['iran '], ['[[scientific reports'], ['bmj global health'], ['bmc evolutionary biology'], [' oxford university press'], ['economic geography'], ['libri ']]",65,12,0,135,0,9,109,0.1906158357771261,0.03519061583577713,0.39589442815249265,0.03519061583577713,0.0,0.26099706744868034,10,"['www.iraqinationality.gov', 'www.cia.gov', 'georgewbush-whitehouse.archives.gov', 'georgewbush-whitehouse.archives.gov', 'www.state.gov', 'www.iraqinationality.gov', 'investpromo.gov', 'www.eia.doe.gov', 'www.eia.doe.gov', 'georgewbush-whitehouse.archives.gov', 'uscis.gov', 'state.gov', 'books.google.com', 'books.google.com', 'www.globalconstructionreview.com', 'www.ft.com', 'www.euromonitor.com', 'abcnews.go.com', 'www.nytimes.com', 'www.youtube.com', 'www.foxnews.com', 'www.bbc.com', 'stadiumdb.com', 'insidearabia.com', 'www.nbcnews.com', 'www.britannica.com', 'www.nytimes.com', 'www.bloomberg.com', 'www.foxnews.com', 'www.lifepersona.com', 'www.theislanderonline.com', 'www.nytimes.com', 'books.google.com', 'www.cnn.com', 'books.google.com', 'www.dangoor.com', 'www.youtube.com', 'foreignpolicy.com', 'www.washingtonpost.com', 'nationalreview.com', 'middleeastvoices.voanews.com', 'www.washingtonpost.com', 'books.google.com', 'www.aljazeera.com', 'www.washingtontimes.com', 'www.foxnews.com', 'www.reuters.com', 'www.bbc.com', 'geography.about.com', 'www.foxnews.com', 'etymonline.com', 'www.huffingtonpost.com', 'edition.cnn.com', 'www.nytimes.com', 'www.jadaliyya.com', 'www.bbc.com', 'dinarprofits.com', 'www.inma-iraq.com', 'www.mnf-iraq.com', 'cnn.com', 'etymonline.com', 'www.reuters.com', 'www.theatlantic.com', 'www.nytimes.com', 'edition.cnn.com', 'america.aljazeera.com', 'www.iraq-businessnews.com', 'asianhistory.about.com', 'www.reuters.com', 'books.google.com', 'iraqinews.com', 'www.nbcnews.com', 'www.britannica.com', 'www.stripes.com', 'www.csmonitor.com', 'usatoday.com', 'books.google.com', 'www.al-monitor.com', 'www.wildlifeextra.com', 'www.cnn.com', 'www.nytimes.com', 'www.thingsasian.com', 'books.google.com', 'www.bartleby.com', 'www.reuters.com', 'www.britannica.com', 'ultrairaq.ultrasawt.com', 'books.google.com', 'www.reuters.com', 'www.aljazeera.com', 'www.newyorker.com', 'www.bbc.com', 'www.business-anti-corruption.com', 'www.arabnews.com', 'www.reuters.com', 'www.aljazeera.com', 'valerieyule.com', 'ca.reuters.com', 'www.reuters.com', 'www.aljazeera.com', 'www.iraqidinar123.com', 'www.france24.com', 'www.aljazeera.com', 'www.sfgate.com', 'articles.latimes.com', 'online.wsj.com', 'www.nytimes.com', 'www.foxnews.com', 'www.arabaviation.com', 'www.reuters.com', 'www.nbcnews.com', 'usatoday30.usatoday.com', 'books.google.com', 'www.washingtonpost.com', 'www.csmonitor.com', 'books.google.com', 'www.alhurra.com', 'www.infoplease.com', 'foreignpolicy.com', 'www.jadaliyya.com', 'waterencyclopedia.com', 'www.nytimes.com', 'books.google.com', 'mertsahinoglu.com', 'www.warprofiteers.com', 'www.reuters.com', 'www.washingtonpost.com', 'www.economist.com', 'www.merriam-webster.com', 'www.reuters.com', 'abcnews.go.com', 'www.britannica.com', 'www.aljazeera.com', 'www.economist.com', 'www.aljazeera.com', 'edition.cnn.com', 'www.reuters.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'www.iraqidinar123.com', 'www.dw.com', 'www.dw.com', 'www.britannica.com', 'www.rfcafe.com', 'edition.cnn.com', 'www.aljazeera.com', 'www.worldhistory.org', 'csis.org', 'www.refworld.org', 'www.irinnews.org', 'sumerian.org', 'domino.un.org', 'www.unicef.org', 'www.internal-displacement.org', 'hrw.org', 'www.iraqicivilsociety.org', '-opcw.org', 'documents1.worldbank.org', 'www.sesrtcic.org', 'www.unesco.org', 'www.climatelinks.org', 'www.longwarjournal.org', 'www.hrw.org', 'stats.oecd.org', 'www.cpa-iraq.org', 'www.worldhistory.org', 'www.unicef.org', 'www.worldhistory.org', 'imf.org', 'www.hrw.org', 'www.sesrtcic.org', 'imf.org', 'www.constituteproject.org', 'data.worldbank.org', 'factcheck.org', 'www.freedomhouse.org', 'www.npr.org', 'domino.un.org', 'medomed.org', 'data2.unhcr.org', 'www.iranicaonline.org', 'www.clingendael.org', 'www.worldhistory.org', 'www.institutkurde.org', 'data.worldbank.org', 'www.imf.org', 'www.genocidewatch.org', 'www.svoboda.org', 'www.cfr.org', 'www.sesrtcic.org', 'www.globalpolicy.org', 'fundforpeace.org', 'www.iraqwatch.org', 'news.un.org', 'www.pewresearch.org', 'rferl.org', 'www.cpa-iraq.org', 'www.constituteproject.org', 'www.unhcr.org', 'www.thenewhumanitarian.org', 'www.opec.org', 'npr.org', 'fundforpeace.org', 'fundforpeace.org', 'ich.unesco.org', 'www.worldhistory.org', 'www.odi.org', 'apps.americanbar.org', 'www.islamopediaonline.org', 'hdr.undp.org', 'whc.unesco.org', ['bioscience'], ['international review of education'], ['intelligence and national security'], ['iran '], ['[[scientific reports'], ['bmj global health'], ['bmc evolutionary biology'], [' oxford university press'], ['economic geography'], ['libri ']]",7515928,Require administrator access (no expiry set),222793,5 May 2001,KoyaanisQatsi ,12311,39,2001-05-05,2001-05,2001
212,212,Sweden,https://en.wikipedia.org/wiki/Sweden,342,6,"['10.1038/s41467-020-19493-3', '10.1093/lawfam/4.2.154', '10.1038/s41561-021-00719-y', None, '10.1175/1520-0493(1900)28[393:tgsm]2.0.co;2', '10.1086/ntj41789232', '33293507', None, None, '11640321', None, None, '7723057', None, None, None, None, None]","[['nature communications'], ['international journal of law'], ['[[nature geoscience'], ['hippokrates. suomen lääketieteen historian seuran vuosikirja'], ['monthly weather review '], ['national tax journal']]",36,10,0,60,0,5,225,0.10526315789473684,0.029239766081871343,0.17543859649122806,0.017543859649122806,0.0,0.15204678362573099,6,"['factfinder.census.gov', 'www.cia.gov', 'www.health.gov', 'www.uspto.gov', 'www.gov', 'www.gov', 'www.gov', 'cia.gov', '2009-2017.state.gov', 'www.cia.gov', 'news.nationalgeographic.com', 'www.nationmaster.com', 'kismeta.com', 'books.google.com', 'www.newstatesman.com', 'books.google.com', 'www.huffingtonpost.com', 'www.economist.com', 'abebooks.com', 'www.nytimes.com', 'www.france24.com', 'books.google.com', 'www.bloomberg.com', 'www.economist.com', 'britannica.com', 'infomotions.com', 'books.google.com', 'www.keepeek.com', 'books.google.com', 'www.nytimes.com', 'query.nytimes.com', 'books.google.com', 'time.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.reuters.com', 'www.economist.com', 'www.americanwest.com', 'dualcitizeninc.com', 'www.bbc.com', 'nationmaster.com', 'www.time.com', 'nationmaster.com', 'www.ferrylines.com', 'books.google.com', 'www.washingtontimes.com', 'www.credit-suisse.com', 'books.google.com', 'www.keepeek.com', 'books.google.com', 'www.keepeek.com', 'concise.britannica.com', 'www.nytimes.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'www.mckinsey.com', 'books.google.com', 'books.google.com', 'query.nytimes.com', 'swedenabroad.com', 'books.google.com', 'www.keepeek.com', 'largestcompanies.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'highbeam.com', 'www.unric.org', 'www.heritage.org', 'www.iclrs.org', 'www.oecd.org', 'www.oecd-ilibrary.org', 'norden.org', 'runeberg.org', 'stats.oecd.org', 'jewishvirtuallibrary.org', 'www.oecd-ilibrary.org', 'pokerfed.org', 'www.imd.org', 'unstats.un.org', 'hdr.undp.org', 'imf.org', 'www.pewresearch.org', 'gtb.ivdnt.org', 'www.sweden.org', 'www.fao.org', 'oecd.org', 'www.childrensfoodtrust.org', 'migrationinformation.org', 'www.iop.org', 'econjwatch.org', 'www.weforum.org', 'www.oecd-ilibrary.org', 'www.oecdbetterlifeindex.org', 'www.un.org', 'hdr.undp.org', 'geographic.org', 'hdr.undp.org', 'www.world-nuclear.org', 'www.globalreligiousfutures.org', 'stats.oecd.org', 'runeberg.org', 'www.oecdbetterlifeindex.org', ['nature communications'], ['international journal of law'], ['[[nature geoscience'], ['hippokrates. suomen lääketieteen historian seuran vuosikirja'], ['monthly weather review '], ['national tax journal']]",5058739,Require administrator access (no expiry set),277914,1 October 2001,DavidSaff ,13440,16,2001-10-01,2001-10,2001
213,213,Norway,https://en.wikipedia.org/wiki/Norway,312,7,"['10.1038/s41467-020-19493-3', None, '10.1016/0048-9697(87)90375-5', '10.1127/0941-2948/2006/0130', '10.1093/biosci/bix014', '10.5194/hess-11-1633-2007', '10.1038/sj.ejhg.5200834', '33293507', '2197762', None, None, '28608869', None, '12173029', '7723057', None, None, None, '5451287', None, None]","[['nature communications'], [' tidsskrift for den norske laegeforening'], ['science of the total environment', 'national academies press'], ['meteorologische zeitschrift'], ['bioscience'], ['hydrology and earth system sciences'], [' european journal of human genetics']]",34,11,0,43,0,1,218,0.10897435897435898,0.035256410256410256,0.13782051282051283,0.022435897435897436,0.0,0.16666666666666666,7,"['2009-2017.state.gov', 'www.cia.gov', 'factfinder.census.gov', 'www.bls.gov', 'www.cia.gov', 'www.bls.gov', 'www.cia.gov', 'factfinder.census.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.usnews.com', 'www.worldbandy.com', 'www.huffingtonpost.com', 'digitaljournal.com', 'www.huffingtonpost.com', 'uk.reuters.com', 'www.embassypages.com', 'www.fifa.com', 'books.google.com', 'www.cnn.com', 'www.britannica.com', '123independenceday.com', 'everyculture.com', 'artcyclopedia.com', 'www.forbes.com', 'www.economist.com', 'books.google.com', 'abcnews.go.com', 'books.google.com', 'dealbook.nytimes.com', 'www.fivb.com', 'forbes.com', 'news.nationalgeographic.com', 'nordictrans.com', 'www.reuters.com', 'encarta.msn.com', 'www.huffingtonpost.com', 'www.ft.com', 'www.economist.com', 'af.reuters.com', 'autoguide.com', 'www.bloomberg.com', 'www.issuesmagazine.com', 'www.britannica.com', 'uk.reuters.com', 'www.lonelyplanet.com', 'hybridcars.com', 'sciencenordic.com', 'www.reuters.com', 'canadianbusiness.com', 'eiu.com', 'norwegianfilm.com', 'religionnews.com', 'climate-data.org', 'www.oecd.org', 'freedomhouse.org', 'norway.org', 'www.weforum.org', 'norway.org', 'norway.org', 'eu-norge.org', 'www.norway.org', 'www.pbs.org', 'www.norway.org', 'www.avere.org', 'norway.org', 'en.rsf.org', 'www.unric.org', 'www.fao.org', 'hdr.undp.org', 'www.oecdbetterlifeindex.org', 'norway.org', 'norway.org', 'panda.org', 'webcitation.org', 'www.transparency.org', 'eplads.norden.org', 'norway.org', 'library.oapen.org', 'www.norway.org', 'www.imf.org', 'hdr.undp.org', 'hdr.undp.org', 'www.galdu.org', 'eoearth.org', 'ourworldindata.org', 'stats.oecd.org', ['nature communications'], [' tidsskrift for den norske laegeforening'], ['science of the total environment', 'national academies press'], ['meteorologische zeitschrift'], ['bioscience'], ['hydrology and earth system sciences'], [' european journal of human genetics']]",21241,Require administrator access (no expiry set),238067,16 November 2001,Eob ,14841,6,2001-11-16,2001-11,2001
214,214,Slavonia,https://en.wikipedia.org/wiki/Slavonia,202,2,"['10.1093/oxfordjournals.ejil.a035834', '10.1136/adc.71.6.540', None, '7726618', None, '1030096']","[['european journal of international law'], [' [[bmj group', ' archives of disease in childhood ']]",4,0,0,50,0,0,146,0.019801980198019802,0.0,0.24752475247524752,0.009900990099009901,0.0,0.0297029702970297,2,"['www.nytimes.com', 'issuu.com', 'books.google.com', 'articles.latimes.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'www.nytimes.com', 'www.nytimes.com', 'www.papukgeopark.com', 'www.vjesnik.com', 'books.google.com', 'www.nytimes.com', 'www.bulgari-istoria-2010.com', 'articles.latimes.com', 'books.google.com', 'www.nytimes.com', 'articles.latimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.encyclopedia.com', 'books.google.com', 'www.nytimes.com', 'www.inyourpocket.com', 'www.vjesnik.com', 'books.google.com', 'books.google.com', 'getbybus.com', 'books.google.com', 'www.kutjevo.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'www.vpz.com', 'books.google.com', 'books.google.com', 'www.duro-dakovic.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'www.nytimes.com', 'h-net.org', 'www.unesco.org', 'www.slobodnaevropa.org', 'hakave.org', ['european journal of international law'], [' [[bmj group', ' archives of disease in childhood ']]",149274,Allow all users (no expiry set),131141,20 November 2002,213.202.122.186 ,855,1,2002-11-20,2002-11,2002
215,215,Bangladesh,https://en.wikipedia.org/wiki/Bangladesh,464,12,"['10.1525/as.1998.38.7.01p0370e', '10.1093/biosci/bix014', '10.1007/bf00175563', '10.1038/sdata.2018.214', '10.1093/heapol/czr025', '10.1017/s0020818318000218', '10.1080/00472337285390641', '10.1186/1475-9276-8-29', '10.1163/156852091x00058', '10.1038/s41467-019-12808-z', '10.1525/as.1972.12.2.01p0190a', '10.1111/j.1467-9272.2005.00494.x', None, '28608869', None, '30375988', '21729917', None, None, '19650938', None, '31664024', None, None, None, '5451287', None, '6207062', None, None, None, '2729304', None, '6820795', None, None]","[['asian survey '], ['bioscience'], ['water'], ['scientific data '], ['health policy and planning '], ['international organization '], ['journal of contemporary asia '], ['international journal for equity in health'], ['journal of the economic and social history of the orient'], ['nature communications'], ['asian survey '], ['the professional geographer ']]",97,36,0,174,0,3,142,0.20905172413793102,0.07758620689655173,0.375,0.02586206896551724,0.0,0.3125,12,"['mof.portal.gov', 'bbs.portal.gov', 'afd.gov', '2009-2017.state.gov', 'ispr.gov', 'bdlaws.minlaw.gov', 'nsc.gov', 'www.mofa.gov', 'www.moef.gov', 'memory.loc.gov', 'bdlaws.minlaw.gov', 'www.btrc.gov', 'ugc.gov', 'state.gov', 'www.bangladesh.gov', 'www.bangladesh.gov', 'www.state.gov', 'afd.gov', '2009-2017.state.gov', 'www.parliament.gov', 'www.bbs.gov', 'visitbangladesh.gov', 'bdlaws.minlaw.gov', 'www.cia.gov', 'ugc.gov', 'dghs.gov', 'mea.gov', 'bdlaws.minlaw.gov', 'www.moedu.gov', 'cia.gov', '2009-2017.state.gov', 'bdlaws.minlaw.gov', '2009-2017.state.gov', 'bdlaws.minlaw.gov', 'www.bangladesh.gov', 'home.treasury.gov', 'bdnews24.com', 'books.google.com', 'books.google.com', 'books.google.com', 'bdchessfed.com', 'books.google.com', 'books.google.com', 'en.prothomalo.com', 'books.google.com', 'books.google.com', 'edition.cnn.com', 'www.dhakatribune.com', 'www.dutchwatersector.com', 'www.dhakatribune.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.youtube.com', 'books.google.com', 'www.youtube.com', 'gulfnews.com', 'books.google.com', 'books.google.com', 'voices.nationalgeographic.com', 'books.google.com', 'archive.dhakatribune.com', 'www.arabnews.com', 'www.daily-sun.com', 'www.diplomat.com', 'www.bbc.com', 'books.google.com', 'global.britannica.com', 'bearprojectbd.weebly.com', 'www.aljazeera.com', 'www.dhakatribune.com', 'archive.dhakatribune.com', 'thediplomat.com', 'books.google.com', 'books.google.com', 'worldpopulationreview.com', 'theodora.com', 'www.bbc.com', 'www.aljazeera.com', 'www.youtube.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'bdnews24.com', 'www.bbc.com', 'www.dw.com', 'www.theatlantic.com', 'cebr.com', 'link.galegroup.com', 'www.aljazeera.com', 'books.google.com', 'books.google.com', 'www.observerbd.com', 'www.youtube.com', 'archive.dhakatribune.com', 'books.google.com', 'opinion.bdnews24.com', 'articles.latimes.com', 'www.britannica.com', 'bdnews24.com', 'academic.eb.com', 'www.financialexpress.com', 'www.dhakatribune.com', 'books.google.com', 'www.photius.com', 'www.britannica.com', 'www.dhakatribune.com', 'www.nationalgeographic.com', 'books.google.com', 'books.google.com', 'www.unb.com', 'books.google.com', 'www.bbc.com', 'google.com', 'bdnews24.com', 'books.google.com', 'www.dailypress.com', 'www.daily-sun.com', 'www.geetabitan.com', 'm.theindependentbd.com', 'books.google.com', 'yourarticlelibrary.com', 'books.google.com', 'thediplomat.com', 'books.google.com', 'www.daily-sun.com', 'theindependentbd.com', 'www.iht.com', 'www.youtube.com', 'sudestada.com', 'books.google.com', 'books.google.com', 'archive.prothom-alo.com', 'cebr.com', 'timesofindia.indiatimes.com', 'books.google.com', 'archive.dhakatribune.com', 'rubaiyat-hossain.com', 'books.google.com', 'govpoliju.com', 'www.dhakatribune.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.britannica.com', 'timesofindia.indiatimes.com', 'www.dhakatribune.com', 'www.dhakachamber.com', 'books.google.com', 'www.economist.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'economictimes.indiatimes.com', 'www.dw.com', 'search.proquest.com', 'books.google.com', 'www.eslteachersboard.com', 'foreignpolicy.com', 'books.google.com', 'www.prothomalo.com', 'www.bbc.com', 'www.discovery.com', 'kantaji.com', 'www.themoscowtimes.com', 'www.reuters.com', 'books.google.com', 'marinelink.com', 'books.google.com', 'bdnes24.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.dhakatribune.com', 'bdnews24.com', 'books.google.com', 'blogs.scientificamerican.com', 'peakbagger.com', 'books.google.com', 'books.google.com', 'books.google.com', 'bdnews24.com', 'www.lonelyplanet.com', 'www.fiercepharmaasia.com', 'books.google.com', 'www.lonelyplanet.com', 'www.youtube.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.aljazeera.com', 'govpoliju.com', 'books.google.com', 'books.google.com', 'www.youtube.com', 'books.google.com', 'www.chevron.com', 'books.google.com', 'news.nationalgeographic.com', 'zeenews.india.com', 'thediplomat.com', 'bdnews24.com', 'www.dhakatribune.com', 'www.dhakatribune.com', 'archive.dhakatribune.com', 'whc.unesco.org', 'www.jstor.org', 'uis.unesco.org', 'www.wssinfo.org', 'bank.org', 'www.worldbank.org', 'www.bangladeshnavy.org', 'en.banglapedia.org', 'www.worldbank.org', 'www.nobelprize.org', 'theismaili.org', 'www.bdhcdelhi.org', 'en.banglapedia.org', 'www.worldbank.org', 'www.futurehealthsystems.org', 'hdr.undp.org', 'www.pewforum.org', 'en.banglapedia.org', 'www.alertnet.org', 'www.wttc.org', 'fao.org', 'www.ti-bangladesh.org', 'www.futurehealthsystems.org', 'en.banglapedia.org', 'freedomhouse.org', 'en.banglapedia.org', 'en.banglapedia.org', 'ilo.org', 'www.wssinfo.org', 'en.banglapedia.org', 'en.banglapedia.org', 'en.banglapedia.org', 'www.iranicaonline.org', 'ejfoundation.org', 'www.amnesty.org', 'en.banglapedia.org', 'persian.packhum.org', 'www.sufismjournal.org', 'lowyinstitute.org', 'treaties.un.org', 'www.imf.org', 'en.banglapedia.org', 'portal.unesco.org', 'www.gwp.org', 'en.banglapedia.org', 'data.worldbank.org', 'features.pewforum.org', 'povertydata.worldbank.org', 'reports.weforum.org', 'www.imf.org', 'en.banglapedia.org', 'freedomhouse.org', 'www.commonwealthofnations.org', 'www.unicef.org', 'www.inm.org', 'en.banglapedia.org', 'www.livelihoods.org', 'data.footprintnetwork.org', 'legal.un.org', 'www.metmuseum.org', 'en.banglapedia.org', 'www.transparency.org', 'www.globalslaveryindex.org', 'www.unesco.org', 'www.iea.org', 'www.bb.org', 'www.amnesty.org', 'www.pewforum.org', 'pewglobal.org', 'www.ti-bangladesh.org', 'www.orfonline.org', 'treaties.un.org', 'www.worldcat.org', 'en.banglapedia.org', 'www.unhcr.org', 'freedomhouse.org', 'web.worldbank.org', 'web.worldbank.org', 'baec.org', 'bti-project.org', 'en.banglapedia.org', 'climatecentral.org', 'carnegieendowment.org', 'constituteproject.org', 'en.banglapedia.org', 'en.banglapedia.org', 'www-wds.worldbank.org', 'www.amnesty.org', 'www.futurehealthsystems.org', 'tonyblairfaithfoundation.org', 'www.asiaticsociety.org', 'en.banglapedia.org', 'www.iranicaonline.org', 'en.banglapedia.org', 'www.nyulawglobal.org', 'www.worldbank.org', 'unesdoc.unesco.org', ['asian survey '], ['bioscience'], ['water'], ['scientific data '], ['health policy and planning '], ['international organization '], ['journal of contemporary asia '], ['international journal for equity in health'], ['journal of the economic and social history of the orient'], ['nature communications'], ['asian survey '], ['the professional geographer ']]",3454,Require administrator access (no expiry set),305911,21 April 2001,Koyaanisqatsi~enwiki ,16932,26,2001-04-21,2001-04,2001
216,216,Offal,https://en.wikipedia.org/wiki/Offal,64,2,"['10.1056/nejme020167', '10.1136/sbmj.0205158', '12540650', None, None, None]","[['new england journal of medicine'], ['student bmj ']]",1,2,0,47,0,0,12,0.015625,0.03125,0.734375,0.03125,0.0,0.078125,2,"['www.foodstandards.gov', 'medlineplus.gov', 'deafnation.com', '973thedawg.com', 'lctabus.com', 'sg.news.yahoo.com', 'naharnet.com', 'kitchendaily.com', 'facts.com', 'www.chilango.com', 'merriam-webster.com', 'www.huffingtonpost.com', 'persianteb.com', 'i57.tinypic.com', 'tribune.com', 'www.usatoday.com', 'www.youtube.com', 'www.youtube.com', 'facts.com', 'travelphotoreport.com', 'foodbycountry.com', 'egyptian-cuisine-recipes.com', 'facts.com', 'uppersia.com', 'facts.com', 'www.bloggang.com', 'www.greenprophet.com', 'digitaljournal.com', 'the-than.com', 'naharnet.com', 'farm1.static.flickr.com', 'bikyamasr.com', 'mawdoo3.com', 'www.nbcnews.com', 'www.klasiktatlar.com', 'chowhound.chow.com', 'books.google.com', 'irishtimes.com', 'christiansofiraq.com', 'www.citylab.com', 'aegis.com', 'books.google.com', 'kale-pache_persianteb.com', 'books.google.com', 'sandandsuccotash.com', 'vagabondish.com', 'washingtonpost.com', 'facts.com', 'www.nytimes.com', 'www.webarchive.org', ['new england journal of medicine'], ['student bmj ']]",342509,Allow all users (no expiry set),79101,16 October 2003,63.80.49.108 ,1415,0,2003-10-16,2003-10,2003
217,217,Culture of Bosnia and Herzegovina,https://en.wikipedia.org/wiki/Culture_of_Bosnia_and_Herzegovina,2,0,[],[],0,0,0,0,0,0,2,0.0,0.0,0.0,0.0,0.0,0.0,0,[],397584,Require autoconfirmed or confirmed access (no expiry set),14583,11 December 2003,212.161.72.152 ,300,0,2003-12-11,2003-12,2003
218,218,Algeria,https://en.wikipedia.org/wiki/Algeria,215,8,"['10.1038/s41467-020-19493-3', '10.1353/cul.2005.0008', '10.1017/s0263718900007810', '10.5944/etfvii.12.1999.2343', '10.1086/423147', '10.1126/science.aau0008', '10.1371/journal.pgen.1002397', '10.3390/resources7030058', '33293507', None, None, None, '15202071', '30498166', '22253600', None, '7723057', None, None, None, '1216069', None, '3257290', None]","[['nature communications'], ['cultural critique'], ['libyan studies'], ['espacio tiempo y forma. serie vii'], ['am. j. hum. genet. '], ['science '], ['plos genetics '], ['resources']]",34,13,0,91,0,1,69,0.15813953488372093,0.06046511627906977,0.4232558139534884,0.037209302325581395,0.0,0.2558139534883721,8,"['www.eia.gov', '2009-2017.state.gov', 'lcweb2.loc.gov', 'www.fco.gov', 'algiers.usembassy.gov', 'www.cia.gov', 'lcweb2.loc.gov', 'cia.gov', 'www.cia.gov', '2009-2017.state.gov', 'www.state.gov', 'webarchive.loc.gov', 'www.cia.gov', 'www.aljazeera.com', 'books.google.com', 'www.lematindalgerie.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.economist.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'khadda.com', 'books.google.com', 'books.google.com', 'www.economist.com', 'www.lebanese-forces.com', 'www.nytimes.com', 'books.google.com', 'books.google.com', 'report.com', 'books.google.com', 'presse-dz.com', 'books.google.com', 'books.google.com', 'articles.cnn.com', 'books.google.com', 'www.upstreamonline.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'african.howzit.msn.com', 'books.google.com', 'www.nytimes.com', 'www.elwatan.com', 'www.upi.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'www1.skysports.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'www.bloomberg.com', 'books.google.com', 'books.google.com', 'www.bbc.com', 'books.google.com', 'magharebia.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'visitwestmanislands.com', 'muslimheritage.com', 'books.google.com', 'algerie-dz.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'tsa-algerie.com', 'books.google.com', 'www.washingtonpost.com', 'books.google.com', 'books.google.com', 'books.google.com', 'fanack.com', 'books.google.com', 'books.google.com', 'www.bbc.com', 'arabicnews.com', 'books.google.com', 'www.zawya.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.frenchpubagency.com', 'books.google.com', 'www.statista.com', 'books.google.com', 'topics.blogs.nytimes.com', 'www.lematindalgerie.com', 'books.google.com', 'www.opec.org', 'www.hrw.org', 'www.unhcr.org', 'www.irinnews.org', 'freedomhouse.org', 'www.unesco.org', 'www.imf.org', 'data.worldbank.org', 'stoneageinstitute.org', 'en.wikisource.org', 'www.freedomhouse.org', 'qantara-med.org', 'whc.unesco.org', 'journals.plos.org', 'www.galtoninstitute.org', 'www.wdl.org', 'archive.ipu.org', 'www.africaneconomicoutlook.org', 'qantara-med.org', 'imf.org', 'hdr.undp.org', 'apn-dz.org', 'worldcat.org', 'rabat.unesco.org', 'nationsonline.org', 'www.globalreligiousfutures.org', 'euromedmonitor.org', 'www.freedomhouse.org', 'www.refugees.org', 'undp-pogar.org', 'www.hrw.org', 'data.footprintnetwork.org', 'www.francophonie.org', 'www.francophonie.org', ['nature communications'], ['cultural critique'], ['libyan studies'], ['espacio tiempo y forma. serie vii'], ['am. j. hum. genet. '], ['science '], ['plos genetics '], ['resources']]",358,Require administrator access (no expiry set),173859,31 October 2001,Corvus13 ,11520,15,2001-10-31,2001-10,2001
219,219,Nigeria,https://en.wikipedia.org/wiki/Nigeria,284,18,"['10.1017/9781108887748', '10.1016/s0048-721x(88)80017-4', '10.1093/oxfordhb/9780198804307.013.13', '10.15177/seefor.14-06', '10.1038/s41467-020-19493-3', '10.4314/jasem.v13i1.55251', None, '10.1016/s0377-8401(99)00131-5', '10.1057/9781137324535', '10.2307/484337', '10.1007/s13644-021-00450-5', '10.1177/002193478101100404', '10.1639/0044-7447(2002)031[0055:wmatfe]2.0.co;2', '10.1111/j.1475-4959.2005.00154.x', '10.4314/as.v8i2.51107', '10.1080/00358535908452221', '10.2752/bewdf/edch1050', '10.2307/1581109', None, None, None, None, '33293507', None, '24739340', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, '7723057', None, '5779393', None, None, None, None, None, None, None, None, None, None, None]","[['cambridge university press'], ['religion '], ['oxford university press'], ['south-east european forestry '], ['nature communications'], ['journal of applied sciences and environmental management'], ['mmwr. morbidity and mortality weekly report'], ['animal feed science and technology'], ['palgrave macmillan'], ['canadian journal of african studies'], [' review of religious research'], ['journal of black studies'], ['ambio'], ['geographical journal'], ['agro-science'], ['[[the round table '], ['berg encyclopedia of world dress and fashion'], ['journal of religion in africa ']]",57,19,0,99,0,8,83,0.2007042253521127,0.06690140845070422,0.3485915492957746,0.06338028169014084,0.0,0.33098591549295775,18,"['files.eric.ed.gov', 'www.fco.gov', 'www.cia.gov', 'www.nigerianstat.gov', 'photos.state.gov', 'nigerianstat.gov', 'www.nigerianstat.gov', 'www.cia.gov', 'www.cia.gov', 'lcweb2.loc.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.fbi.gov', 'www.cia.gov', 'www.cia.gov', 'www.state.gov', 'www.cia.gov', 'www.time.com', 'www.nigerdeltacongress.com', 'www.nationsencyclopedia.com', 'www.onlinenigeria.com', 'www.channelstv.com', 'myondostate.com', 'www.nytimes.com', 'www.tribune.com', 'www.csmonitor.com', 'books.google.com', 'www.nytimes.com', 'www.vanguardngr.com', 'www.cnn.com', 'www.zambianwatchdog.com', 'www.mydailynewswatchng.com', 'books.google.com', 'www.economist.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.vanguardngr.com', 'books.google.com', 'www.si.com', 'books.google.com', 'www.cgwic.com', 'africa.com', 'www.fivb.com', 'books.google.com', 'www.reuters.com', 'hautefashionafrica.com', 'www.bellanaija.com', 'pacmar.com', 'www.csmonitor.com', 'books.google.com', 'www.cnbc.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'www.vanguardngr.com', 'www.theatlantic.com', 'www.sunnewsonline.com', 'books.google.com', 'www.economist.com', 'www.msn.com', 'books.google.com', 'www.africanews.com', 'africabasket.com', 'books.google.com', 'litencyc.com', 'books.google.com', 'www.thestandard.com', 'www.thearda.com', 'www.reuters.com', 'america.aljazeera.com', 'www.innosonvehicles.com', 'fiba.com', 'books.google.com', 'www.thehistoryville.com', 'www.thisdaylive.com', 'books.google.com', 'www.sunnewsonline.com', 'www.bbc.com', 'www.nigeriasun.com', 'www.punchng.com', 'www.ethnologue.com', 'www.bbc.com', 'www.ethnologue.com', 'www.thisdaylive.com', 'www.economist.com', 'www.newframe.com', 'edition.cnn.com', 'books.google.com', 'www.punchng.com', 'books.google.com', 'naijalitz.com', 'www.vanguardngr.com', 'rainforests.mongabay.com', 'www.forbes.com', 'books.google.com', 'africanspotlight.com', 'africafootunited.com', 'encarta.msn.com', 'af.reuters.com', 'www.vanguardngr.com', 'allafrica.com', 'books.google.com', 'www.thenigerianvoice.com', 'afp.google.com', 'www.economist.com', 'www.vanguardngr.com', 'www.cgwic.com', 'news.mongabay.com', 'www.washingtonpost.com', 'news2.onlinenigeria.com', 'etymonline.com', 'books.google.com', 'www.worldcat.org', 'www.refworld.org', 'freedomhouse.org', 'www.casade.org', 'www.nigeria-law.org', 'features.pewforum.org', 'www.prb.org', 'profiles.countdown2030.org', 'worldcurling.org', 'hdr.undp.org', 'treaties.un.org', 'www.pewglobal.org', 'hdr.undp.org', 'wwrn.org', 'wwrn.org', 'www.cgdev.org', 'www.africaleadership.org', 'www.pewresearch.org', 'esa.un.org', 'www.pewforum.org', 'www.assatashakur.org', 'www.npr.org', 'hdr.undp.org', 'www.cambridge.org', 'www.efccnigeria.org', 'www.imf.org', 'metmuseum.org', 'features.pewforum.org', 'www.americamagazine.org', 'pewforum.org', 'heapol.oxfordjournals.org', 'www.africa-union.org', 'wiwavshell.org', 'www.nti.org', 'www.un.org', 'www.bahai.org', 'www.ohchr.org', 'pewforum.org', 'www.cfr.org', 'www.pewresearch.org', 'www.radionetherlandsarchives.org', 'hdr.undp.org', 'iea.org', 'nasarawastate.org', 'www.worldbank.org', 'www.efccnigeria.org', 'yorubanation.org', 'www.alertnet.org', 'www.iucngisd.org', 'www.cambridge.org', 'www.eueom-ng.org', 'data.worldbank.org', 'worldcat.org', 'www.migrationinformation.org', 'www.pbs.org', 'data.worldbank.org', 'www.eldis.org', ['cambridge university press'], ['religion '], ['oxford university press'], ['south-east european forestry '], ['nature communications'], ['journal of applied sciences and environmental management'], ['mmwr. morbidity and mortality weekly report'], ['animal feed science and technology'], ['palgrave macmillan'], ['canadian journal of african studies'], [' review of religious research'], ['journal of black studies'], ['ambio'], ['geographical journal'], ['agro-science'], ['[[the round table '], ['berg encyclopedia of world dress and fashion'], ['journal of religion in africa ']]",21383,Require administrator access (no expiry set),206407,25 May 2001,KoyaanisQatsi ,9356,26,2001-05-25,2001-05,2001
220,220,Ethiopia,https://en.wikipedia.org/wiki/Ethiopia,475,29,"['10.1525/ae.1975.2.4.02a00030', '10.1038/nature03258', '10.1038/news050214-10', '10.1126/science.aaw8942', '10.1186/s13033-017-0144-4', '10.1126/science.1153717', '10.1016/j.jhevol.2017.04.004', '10.1093/aob/mcy214', '10.1038/nature.2017.22114', '10.1038/s41467-020-19493-3', '10.1371/journal.pone.0216716', '10.1371/journal.pone.0078092', '10.1017/s0022278x00055233', '10.1038/nature01669', '10.3406/galim.2012.1993', '10.1017/s0041977x00056731', '10.1098/rspb.2016.0792', '10.4314/ahs.v17i3.9', '10.2307/1357309', '10.1126/science.1078208', '10.2307/216612', '10.1016/0169-5150(91)90022-d', '10.1080/23311932.2019.1613770', '10.1093/jhmas/xxi.2.95', '10.1080/01436599814415', '10.1017/s0041977x00144209', '10.1098/rspb.1976.0061', None, '15716951', None, '31395781', '28603550', '18292342', '28552208', '30715125', None, '33293507', '31071181', '24236011', None, '12802332', None, None, None, '29085394', None, '12714734', None, None, None, '5326887', None, None, '11482', None, None, None, None, '5465569', None, None, '6526316', None, '7723057', '6508696', '3827237', None, None, None, None, '4920324', '5656212', None, None, None, None, None, None, None, None, None]","[[' american ethnologist'], [' nature '], ['[[nature '], ['science'], ['international journal of mental health systems'], ['[[science '], ['journal of human evolution'], ['annals of botany'], ['[[nature '], ['nature communications'], ['plos one'], ['plos one '], ['the journal of modern african studies '], [' nature'], ['gazette du livre médiéval'], ['bulletin of the school of oriental and african studies '], ['proc. r. soc. b'], ['african health sciences '], ['bulletin of the american schools of oriental research '], [' science '], ['international journal of african studies '], [' agricultural economics'], ['cogent food '], [' journal of the history of medicine and allied sciences'], ['third world quarterly '], [' bulletin of the school of oriental and african studies'], ['proceedings of the royal society of london. series b. biological sciences']]",78,25,0,186,0,7,152,0.16421052631578947,0.05263157894736842,0.391578947368421,0.061052631578947365,0.0,0.27789473684210525,27,"['www.cia.gov', 'www.csa.gov', 'www.csa.gov', 'memory.loc.gov', 'www.cia.gov', 'memory.loc.gov', 'www.ethiopia.gov', '2009-2017.state.gov', 'www.cia.gov', 'www.ethiopia.gov', 'www.csa.gov', 'dait.interno.gov', 'www.cia.gov', 'www.ena.gov', '2009-2017.state.gov', 'www.csa.gov', 'www.csa.gov', 'www.ethiopia.gov', 'cia.gov', 'www.ethiopia.gov', 'www.csa.gov', 'www.cia.gov', 'www.mwud.gov', 'www.fsc.gov', 'memory.loc.gov', 'nationalgeographic.com', 'allaboutethio.com', 'www.styaredcuisine.com', 'www.ethiopianreporter.com', 'www.nytimes.com', 'books.google.com', 'www.france24.com', 'rainforests.mongabay.com', 'www.aa.com', 'books.google.com', 'books.google.com', 'www.reuters.com', 'www.africanews.com', 'www.bbc.com', 'www.bloomberg.com', 'books.google.com', 'www.google.com', 'www.hydroworld.com', 'www.smithsonianmag.com', 'www.nytimes.com', 'www.theglobeandmail.com', 'af.reuters.com', 'www.africaw.com', 'books.google.com', 'books.google.com', 'www.cnn.com', 'books.google.com', 'allaboutethio.com', 'books.google.com', 'railwaygazette.com', 'www.tigraionline.com', 'tusker.com', 'www.ethiopia-insight.com', 'www.africanews.com', 'www.bbc.com', 'apnews.com', 'worldpopulationreview.com', 'w7news.com', 'www.youtube.com', 'qz.com', 'books.google.com', 'books.google.com', 'www.bbc.com', 'railwaygazette.com', 'www.aljazeera.com', 'www.nature.com', 'www.bbc.com', 'books.google.com', 'gizmodo.com', 'www.startribune.com', 'www.africanews.com', 'www.ethiopianairlines.com', 'wendybelcher.com', 'www.reuters.com', 'infomineo.com', 'www.nazret.com', 'www.news24.com', 'apnews.com', 'www.google.com', 'books.google.com', 'cyberethiopia.com', 'books.google.com', 'www.time.com', 'www.reuters.com', 'www.google.com', 'books.google.com', 'www.upi.com', 'www.aljazeera.com', 'www.bbc.com', 'www.washingtonpost.com', 'www.newsweek.com', 'vislardica.com', 'terradaily.com', 'books.google.com', 'www.usatoday.com', 'english.people.com', 'www.bbc.com', 'addisstandard.com', 'www.aljazeera.com', 'www.thespruceeats.com', 'www.washingtonpost.com', 'rainforests.mongabay.com', 'newbusinessethiopia.com', 'www.youtube.com', 'www.somtribune.com', 'www.bbc.com', 'www.time.com', 'highbeam.com', 'www.ym.com', 'www.britannica.com', 'www.re-thinkingthefuture.com', 'www.nytimes.com', 'www.ethiopia-insight.com', 'livescience.com', 'www.re-thinkingthefuture.com', 'books.google.com', 'www.newsweek.com', 'www.ethnologue.com', 'www.internetlivestats.com', 'www.miceethiopia.com', 'www.nytimes.com', 'books.google.com', 'www.bbc.com', 'realitysandwich.com', 'arstechnica.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'www.economist.com', 'www.smithsonianmag.com', 'www.ethiopianairlines.com', 'books.google.com', 'www.cattlenetwork.com', 'www.reuters.com', 'www.aljazeera.com', 'www.africanews.com', 'www.france24.com', 'books.google.com', 'books.google.com', 'www.dailystar.com', 'www.reuters.com', 'www.google.com', 'books.google.com', 'www.bbc.com', 'allafrica.com', 'www.google.com', 'www.ezega.com', 'www.ethiopiaobserver.com', 'www.washingtonpost.com', 'www.africanews.com', 'www.newsweek.com', 'www.civicwebs.com', 'graphics.eiu.com', 'www.dailysabah.com', 'www.time.com', 'www.bbc.com', 'edition.cnn.com', 'www.nytimes.com', 'www.nationsencyclopedia.com', 'books.google.com', 'www.cattlenetwork.com', 'www.youtube.com', 'photius.com', 'www.horndaily.com', 'www.aljazeera.com', 'books.google.com', 'airport-authority.com', 'endageredspecie.com', 'ethiopianreporter.com', 'ladywriteronline.wordpress.com', 'www.voanews.com', 'eduplace.com', 'www.aljazeera.com', 'books.google.com', 'www.biblegateway.com', 'www.bbc.com', 'www.aljazeera.com', 'www.google.com', 'www.aljazeera.com', 'aljazeera.com', 'ethiopianhistory.com', 'addistribune.com', 'www.rollingstone.com', 'www.business-anti-corruption.com', 'www.nytimes.com', 'www.nytimes.com', 'www.britannica.com', 'aljazeera.com', 'venturesafrica.com', 'www.reuters.com', 'reuters.com', 'allafrica.com', 'akhrailway.com', 'irinnews.com', 'edition.cnn.com', 'www.boundless.com', 'www.biblegateway.com', 'www.tadias.com', 'cnn.com', 'www.bbc.com', 'books.google.com', 'www.washingtonpost.com', 'www.kilil5.com', 'allaboutethio.com', 'qz.com', 'www.time.com', 'www.worldbank.org', 'www.irinnews.org', 'data.uis.unesco.org', 'prb.org', 'www.amnesty.org', 'www.et.undp.org', 'www.irinnews.org', 'www.refugees.org', 'whc.unesco.org', 'freedomhouse.org', 'www.olympic.org', 'www.hrw.org', 'www.etharc.org', 'www.olympic.org', 'www.healthdata.org', 'www.imf.org', 'blackpast.org', 'www.hrw.org', 'www.wateraid.org', 'www.worldcat.org', 'pewglobal.org', 'www.nationalgeographic.org', 'planipolis.iiep.unesco.org', 'data.worldbank.org', 'hrw.org', 'worldbank.org', 'www.dskmariam.org', 'www.freedomhouse.org', 'ooni.torproject.org', 'imf.org', 'npr.org', 'www.africanculturalcenter.org', 'data.un.org', 'britishmuseum.org', 'unesdoc.unesco.org', 'www.khanacademy.org', 'www.worldbank.org', 'www.africa-eu-partnership.org', 'www.ilo.org', 'worldcat.org', 'avibase.bsc-eoc.org', 'www.weforum.org', 'data.worldbank.org', 'www.imf.org', 'www.wilsoncenter.org', 'data.worldbank.org', 'totalitarismo.altervista.org', 'www.worldhistory.org', 'www.worldbank.org', 'www.amnesty.org', 'www.jstor.org', 'npr.org', 'hdr.undp.org', 'www.worldbank.org', 'ethnomed.org', 'oaklandinstitute.org', 'worldbank.org', 'ethiopia.un.org', 'gargaaraoromopc.org', 'developmentprogress.org', 'www.odi.org', 'www.worldbank.org', 'rightlivelihood.org', 'mdgs.un.org', 'freedomhouse.org', 'hdr.undp.org', 'www.irinnews.org', 'www.worldhistory.org', 'kolibri.teacherinabox.org', 'jewishvirtuallibrary.org', 'www.npr.org', 'www.oaklandinstitute.org', 'www.worldcat.org', 'www.hrw.org', 'trialinternational.org', 'trialinternational.org', 'unicef.org', 'www.animalinfo.org', [' american ethnologist'], [' nature '], ['[[nature '], ['science'], ['international journal of mental health systems'], ['[[science '], ['journal of human evolution'], ['annals of botany'], ['[[nature '], ['nature communications'], ['plos one'], ['plos one '], ['the journal of modern african studies '], [' nature'], ['gazette du livre médiéval'], ['bulletin of the school of oriental and african studies '], ['proc. r. soc. b'], ['african health sciences '], ['bulletin of the american schools of oriental research '], [' science '], ['international journal of african studies '], [' agricultural economics'], ['cogent food '], [' journal of the history of medicine and allied sciences'], ['third world quarterly '], [' bulletin of the school of oriental and african studies'], ['proceedings of the royal society of london. series b. biological sciences']]",187749,Require administrator access (no expiry set),297790,30 September 2001,Ap ,17212,84,2001-09-30,2001-09,2001
221,221,Iceland,https://en.wikipedia.org/wiki/Iceland,307,8,"['10.1073/pnas.0902522107', '10.2307/2173366', '10.1093/petrology/5.3.435', '10.1016/s0360-3199(99)00077-4', '10.1111/0021-8294.00054', '10.5194/acpd-3-1599-2003', '10.1001/archsurg.141.2.199', '10.1086/303046', '20212157', '11630504', None, None, None, None, '16490899', '10931763', '2851789', None, None, None, None, None, None, '1287529']","[['proceedings of the national academy of sciences '], ['population studies '], ['journal of petrology '], ['international journal of hydrogen energy '], ['journal for the scientific study of religion '], ['atmospheric chemistry and physics discussions '], [' arch surg'], [' american journal of human genetics']]",43,9,0,61,0,4,182,0.14006514657980457,0.029315960912052116,0.1986970684039088,0.026058631921824105,0.0,0.19543973941368079,8,"['www.cia.gov', 'cia.gov', 'www.cia.gov', 'www.gov', 'www.gov', 'www.gov', 'www.gov', 'state.gov', 'factfinder.census.gov', 'www.bloomberg.com', 'api.nationalgeographic.com', 'www.icelandreview.com', 'www.huffingtonpost.com', 'books.google.com', 'books.google.com', 'www.eiu.com', 'www.visiticeland.com', 'nasdaqomx.com', 'www.wingia.com', 'fortune.com', 'dualcitizeninc.com', 'rottentomatoes.com', 'www.nytimes.com', 'www.icelandreview.com', 'www.bbc.com', 'www.thedailybeast.com', 'kefairport.com', 'www.mensjournal.com', 'www.reuters.com', 'books.google.com', 'blogs.indiewire.com', 'www.nytimes.com', 'www.thehistoryofcanadapodcast.com', 'books.google.com', 'artsbeat.blogs.nytimes.com', 'www.vanityfair.com', 'findarticles.com', 'www.icelandicroots.com', 'uk.reuters.com', 'guinnessworldrecords.com', 'www.travelade.com', 'news.nationalgeographic.com', 'www.usatoday.com', 'www.thehistoryofcanadapodcast.com', 'www.icelandreview.com', 'books.google.com', 'goscandinavia.about.com', 'icelandreview.com', 'guinnessworldrecords.com', 'edition.cnn.com', 'www.bbc.com', 'www.washingtontimes.com', 'www.france24.com', 'www.icelandicroots.com', 'www.biography.com', 'travel-wonders.com', 'ngm.nationalgeographic.com', 'www.iht.com', 'edition.cnn.com', 'www.guinnessworldrecords.com', 'www.engadget.com', 'askjaenergy.com', 'www.guinnessworldrecords.com', 'www.worldatlas.com', 'www.nytimes.com', 'edition.cnn.com', 'nationmaster.com', 'dannyreviews.com', 'www.rigzone.com', 'books.google.com', 'askjaenergy.org', 'www.freedomhouse.org', 'www.imf.org', 'oecd.org', 'oecd.org', 'www.norden.org', 'unesdoc.unesco.org', 'oecd.org', 'voxeu.org', 'www.askjaenergy.org', 'oecd.org', 'archaeology.org', 'worldenergy.org', 'www.visionofhumanity.org', 'www.ilo.org', 'hdr.undp.org', 'ipu.org', 'www.un.org', 'www.chabad.org', 'oecd.org', 'stats.oecd.org', 'oecd.org', 'www3.weforum.org', 'iceland.org', 'oecdbetterlifeindex.org', 'oscars.org', 'members.weforum.org', 'members.weforum.org', 'www.nordicenergysolutions.org', 'esa.un.org', 'npr.org', 'heritage.org', 'stats.oecd.org', 'askjaenergy.org', 'hdr.undp.org', 'oecdbetterlifeindex.org', 'www.heritage.org', 'www.globalinnovationindex.org', 'askjaenergy.org', 'hdr.undp.org', 'hdr.undp.org', 'cpi.transparency.org', 'oecd.org', ['proceedings of the national academy of sciences '], ['population studies '], ['journal of petrology '], ['international journal of hydrogen energy '], ['journal for the scientific study of religion '], ['atmospheric chemistry and physics discussions '], [' arch surg'], [' american journal of human genetics']]",14531,Require administrator access (no expiry set),193474,3 August 2001,Pinkunicorn ,11408,2,2001-08-03,2001-08,2001
222,222,Belgium,https://en.wikipedia.org/wiki/Belgium,278,9,"['10.1159/000013462', '10.4000/etudesrurales.9499', '10.1093/biosci/bix014', '10.1038/s41467-020-19493-3', '10.3406/rbph.1925.6335', '10.1080/01434630208666453', '10.5194/hess-11-1633-2007', '10.3390/resources7030058', '10.2307/3711670', '10213829', None, '28608869', '33293507', None, None, None, None, None, None, None, '5451287', '7723057', None, None, None, None, None]","[['american journal of nephrology'], [' études rurales '], ['bioscience'], ['nature communications'], ['revue belge de philologie et d'], ['journal of multilingual and multicultural development '], ['[[hydrology and earth system sciences'], ['resources'], [' sociological analysis ']]",37,10,0,66,0,1,157,0.13309352517985612,0.03597122302158273,0.23741007194244604,0.03237410071942446,0.0,0.2014388489208633,9,"['nces.ed.gov', '2009-2017.state.gov', 'www.cia.gov', '2009-2017.state.gov', 'www.cia.gov', 'www.cia.gov', 'belgium.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.france24.com', 'books.google.com', 'www.epicurious.com', 'uk.encarta.msn.com', 'www.senses-artnouveau.com', 'blogs.wsj.com', 'wwar.com', 'www.questia.com', 'www.globalpost.com', 'www.cnn.com', 'www.france24.com', 'uk.encarta.msn.com', 'www.euractiv.com', 'edit.britannica.com', 'www.authorama.com', 'www.fifa.com', 'www.britannica.com', 'foodproductiondaily.com', 'wwar.com', 'www.questia.com', 'www.belgianexperts.com', '(alibris.com', 'www.epicurious.com', 'uk.encarta.msn.com', 'www.expatica.com', 'dw.com', 'houbi.com', 'www.visitbelgium.com', 'articles.chicagotribune.com', 'www.inbev.com', 'www.ft.com', 'books.google.com', 'books.google.com', 'www.numbeo.com', 'books.google.com', 'www.globalgourmet.com', 'www.fifa.com', 'dw.com', 'www.ethnologue.com', 'www.france24.com', 'books.google.com', 'books.google.com', 'www.senses-artnouveau.com', 'www.ethnologue.com', 'nytimes.com', 'www.britannica.com', 'www.xpats.com', 'www.expatica.com', 'books.google.com', 'cnn.com', 'www.globalgourmet.com', 'www.eubusiness.com', 'www.123independenceday.com', 'www1.uol.com', 'cnn.com', 'wwar.com', 'www.reuters.com', 'fashionworlds.blogspot.com', 'www.sfgate.com', 'www.belgianexperts.com', 'wwar.com', 'www.portofantwerp.com', 'www.authorama.com', 'sites.google.com', 'www.filmbirth.com', 'www.filmbirth.com', 'www.constituteproject.org', 'nobelprize.org', 'journals.openedition.org', 'iso.org', 'hdr.undp.org', 'www.oecd.org', 'www.ncata.org', 'electionresources.org', 'www.imf.org', 'www.fromoldbooks.org', 'ourworldindata.org', 'whc.unesco.org', 'www.metmuseum.org', 'kp.org', 'hdr.undp.org', 'www.amnh.org', 'www.britishcouncil.org', 'whc.unesco.org', 'zacat.gesis.org', 'www.metmuseum.org', 'www.bh.org', 'hdr.undp.org', 'undp.org', 'zacat.gesis.org', 'www.fromoldbooks.org', 'www.unrisd.org', 'www.ncata.org', 'www.wsws.org', 'hdr.undp.org', 'whc.unesco.org', 'stats.oecd.org', 'www.metmuseum.org', 'www.britishcouncil.org', 'www.catholiceducation.org', 'www.oecd.org', 'data.footprintnetwork.org', 'www.unesco.org', ['american journal of nephrology'], [' études rurales '], ['bioscience'], ['nature communications'], ['revue belge de philologie et d'], ['journal of multilingual and multicultural development '], ['[[hydrology and earth system sciences'], ['resources'], [' sociological analysis ']]",3343,Require administrator access (no expiry set),204197,27 October 2001,PaulFontaine ,11526,12,2001-10-27,2001-10,2001
223,223,Circassians,https://en.wikipedia.org/wiki/Circassians,201,7,"['10.1017/s0020743817000617', '10.1111/j.1467-6443.2005.00262.x', 'abs/10.1080/13537110701293500', '10.1016/j.lingua.2003.06.003', '10.1093/acprof:oso/9780195177756.001.0001', '10.1163/1573384054068123', '10.1126/science.1153717', None, None, None, None, None, None, '18292342', None, None, None, None, None, None, None]","[['international journal of middle east studies'], ['journal of historical sociology'], ['nationalism and ethnic politics '], ['lingua'], ['oxford university press'], ['iran and the caucasus'], ['science']]",27,7,0,46,0,0,114,0.13432835820895522,0.03482587064676617,0.22885572139303484,0.03482587064676617,0.0,0.20398009950248755,7,"['2001.ukrcensus.gov', '2001.ukrcensus.gov', 'memory.loc.gov', '2001.ukrcensus.gov', 'belstat.gov', '2001.ukrcensus.gov', 'www.toplukatalog.gov', 'books.google.com', 'jinepsgazetesi.com', 'www.al-monitor.com', 'www.nytimes.com', 'circassianworld.com', 'books.google.com', 'circassianworld.blogspot.com', 'books.google.com', 'forward.com', 'www.echoesfromjordan.com', 'books.google.com', 'books.google.com', 'books.google.com', 'world.time.com', 'www.nytimes.com', 'books.google.com', 'www.youtube.com', 'books.google.com', 'books.google.com', 'www.trtworld.com', 'www.circassianworld.com', 'i-cias.com', 'www.circassianworld.com', 'www.internethaber.com', 'books.google.com', 'www.youtube.com', 'www.circassianworld.com', 'books.google.com', 'www.myjewishlearning.com', 'books.google.com', 'books.google.com', 'archive.constantcontact.com', 'books.google.com', 'books.google.com', 'caucasustimes.com', 'www.circassianworld.com', 'abkhazworld.com', 'www.reuters.com', 'youtube.com', 'www.britannica.com', 'books.google.com', 'www.circassiancenter.com', 'www.britannica.com', 'books.google.com', 'www.circassianworld.com', 'books.google.com', 'elalliance.org', 'bianet.org', 'www.iranicaonline.org', 'www.iranicaonline.org', 'worldcat.org', 'minorityrights.org', 'www.aheku.org', 'kafkas.org', 'minorityrights.org', 'sreda.org', 'www.iranicaonline.org', 'en.wikipedia.org', 'jamestown.org', 'www.iranicaonline.org', 'www.jamestown.org', 'www.cerkesya.org', 'sreda.org', 'www.jamestown.org', 'www.rferl.org', 'www.orsam.org', 'weekly.ahram.org', 'www.jewishvirtuallibrary.org', 'minorityrights.org', 'sreda.org', 'russiaprofile.org', 'www.ponarseurasia.org', 'www.jamestown.org', ['international journal of middle east studies'], ['journal of historical sociology'], ['nationalism and ethnic politics '], ['lingua'], ['oxford university press'], ['iran and the caucasus'], ['science']]",517916,Allow all users (no expiry set),130297,10 March 2004,ChrisO~enwiki ,2735,15,2004-03-10,2004-03,2004
224,224,Hamburg,https://en.wikipedia.org/wiki/Hamburg,170,0,[],[],11,1,0,30,0,0,129,0.06470588235294118,0.0058823529411764705,0.17647058823529413,0.0,0.0,0.07058823529411765,0,"['ftp.atdd.noaa.gov', 'de.statista.com', 'www.weather-atlas.com', 'www.weatherbase.com', 'de.statista.com', 'hinduonnet.com', 'gl-bfg.com', 'europeupclose.com', 'gl-bfg.com', 'www.boosey.com', 'news.bloodhorse.com', 'hinduonnet.com', 'ning.com', 'soccerlens.com', 'aapa.files.cms-plus.com', 'www.reeperbahnfestival.com', 'kartenseite.files.wordpress.com', 'de.statista.com', 'www.outsports.com', 'mercer.com', 'www.handelsblatt.com', 'hamburgwarriors.com', 'moovitapp.com', 'moovitapp.com', 'www.usatoday.com', 'discogs.com', 'www.airbus.com', 'movielocations.com', 'archnewsnow.com', 'travel-library.com', 'www.merriam-webster.com', 'www.iaaf.org', 'www.audubonmagazine.org', 'hdi.globaldatalab.org', 'en.wtcf.org', 'aapa-ports.org', 'www.sidmartinbio.org', 'www.iaaf.org', 'www.awchamburg.org', 'chabad.org', 'freimaurer.org', 'kreativgesellschaft.org']",13467,Allow all users (no expiry set),141398,13 November 2001,H.J. ,5434,5,2001-11-13,2001-11,2001
225,225,Maharashtra,https://en.wikipedia.org/wiki/Maharashtra,322,7,"['10.1353/jod.2005.0018', '10.4103/0975-2870.118294', '10.1007/s12040-013-0294-y', '10.1080/00220380802265108', '10.1109/igarss.2017.8128250', None, None, None, None, None, None, None, None, None, None]","[['journal of democracy '], ['medical journal of dr. d.y. patil university '], ['journal of earth system science '], ['the journal of development studies '], ['ieee international geoscience and remote sensing symposium ']]",31,45,0,147,0,0,92,0.09627329192546584,0.13975155279503104,0.45652173913043476,0.021739130434782608,0.0,0.2577639751552795,5,"['www.maharashtratourism.gov', 'farmech.gov', 'censusindia.gov', 'maharashtrabiodiversityboard.gov', 'cad.gujarat.gov', 'msrtc.gov', 'mmrda.maharashtra.gov', 'www.maharashtratourism.gov', 'www.maharashtra.gov', 'www.cr.indianrailways.gov', 'www.maha-arogya.gov', 'tourism.gov', 'www.maha-arogya.gov', 'www.censusindia.gov', 'mahades.maharashtra.gov', 'www.kolhapurcorporation.gov', 'mpcb.gov', 'www.maharashtra.gov', 'censusindia.gov', 'maharashtratourism.gov', 'www.dipp.gov', 'pibmumbai.gov', 'knowindia.gov', 'www.wr.indianrailways.gov', 'nrhm.gov', 'www.mahapanchayat.gov', 'www.maharashtra.gov', 'www.maharashtratourism.gov', 'www.censusindia.gov', 'mahades.maharashtra.gov', 'www.maharashtra.gov', 'mahades.maharashtra.gov', 'www.censusindia.gov', 'mpcb.gov', 'maharashtratourism.gov', 'censusindia.gov', 'www.maharashtra.gov', 'maha.gov', 'ffo.gov', 'arogya.maharashtra.gov', 'www.mpcb.gov', 'pdf.usaid.gov', 'maharashtrabiodiversityboard.gov', 'censusindia.gov', 'krishi.maharashtra.gov', 'books.google.com', 'books.google.com', 'books.google.com', 'www.mahasec.com', 'www.amazingmaharashtra.com', 'books.google.com', 'economictimes.indiatimes.com', 'books.google.com', 'www.thehindu.com', 'www.frontierweekly.com', 'www.educationinfoindia.com', 'articles.economictimes.indiatimes.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.atptour.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'rediff.com', 'greencleanguide.com', 'books.google.com', 'www.maharashtrastat.com', 'books.google.com', 'rediff.com', 'books.google.com', 'marathiheritage.com', 'books.google.com', 'cities.expressindia.com', 'www.firstpost.com', 'm.timesofindia.com', 'www.thehindubusinessline.com', 'books.google.com', 'www.discoveredindia.com', 'www.economist.com', 'www.fifaworldcuphub.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.pppinindia.com', 'archive.indianexpress.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.espncricinfo.com', 'www.populationindia.com', 'books.google.com', 'books.google.com', 'exchange4media.com', 'www.maharashtrastat.com', 'www.marathiheritage.com', 'timesofindia.indiatimes.com', 'discoveredindia.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'thehindu.com', 'books.google.com', 'www.jagran.com', 'm.divyamarathi.bhaskar.com', 'delhimumbaiindustrialcorridor.com', 'www.dnaindia.com', 'www.financialexpress.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'indianpowersector.com', 'm.timesofindia.com', 'timesofindia.indiatimes.com', 'centralclusteruupgs.wordpress.com', 'www.eflifans.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'www.veethi.com', 'www.discoveredindia.com', 'archive.indianexpress.com', 'www.amarujala.com', 'rwitc.com', 'books.google.com', 'books.google.com', 'www.efli.com', 'books.google.com', 'books.google.com', 'www.deccanchronicle.com', 'www.espncricinfo.com', 'www.mumbaicricket.com', 'timesofindia.indiatimes.com', 'www.firstpost.com', 'www.tabletmag.com', 'indianexpress.com', 'maharashtracongress.com', 'rjelal.com', 'books.google.com', 'books.google.com', 'www.financialexpress.com', 'timesofindia.indiatimes.com', 'ehealth.eletsonline.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.dailypioneer.com', 'www.esakal.com', 'indianexpress.com', 'zeenews.india.com', 'books.google.com', 'marathiheritage.com', 'www.hindustantimes.com', 'www.mahammb.com', 'www.shvoong.com', 'www.britannica.com', 'www.hindustantimes.com', 'books.google.com', 'm.timesofindia.com', 'www.hindustantimes.com', 'books.google.com', 'books.google.com', 'www.rediff.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.shvoong.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'content.time.com', 'rwitc.com', 'www.thehindubusinessline.com', 'indiatimes.com', 'food.ndtv.com', 'indianexpress.com', 'books.google.com', 'books.google.com', 'books.google.com', 'archive.tehelka.com', 'timesofindia.indiatimes.com', 'www.proquest.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.maharashtraopen.com', 'discoveredindia.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.oocities.org', 'countercurrents.org', 'www-cambridge-org.wikipedialibrary.idm.oclc.org', 'www.unicef.org', 'linguistlist.org', 'www.jstor.org', 'www.coep.org', 'mercindia.org', 'csi-sigegov.org', 'electricitygovernance.wri.org', 'www.in.undp.org', 'www.cehat.org', 'www.auditbureau.org', 'www.in.undp.org', 'karmayog.org', 'aicte-india.org', 'globaldatalab.org', 'ibef.org', 'www.ccmaharashtra.org', 'www.mssidc.org', 'www.auditbureau.org', 'ncte-india.org', 'www.madcindia.org', 'www.jstor.org', 'www.rbi.org', 'sikhinstitute.org', 'lawsofindia.org', 'mcaer.org', 'www.rbi.org', 'rbi.org', 'www.indiapress.org', ['journal of democracy '], ['medical journal of dr. d.y. patil university '], ['journal of earth system science '], ['the journal of development studies '], ['ieee international geoscience and remote sensing symposium ']]",20629,"Require autoconfirmed or confirmed access (08:20, 25 February 2023)",217469,1 December 2001,128.101.45.xxx ,9079,95,2001-12-01,2001-12,2001
226,226,Kazakhstan,https://en.wikipedia.org/wiki/Kazakhstan,291,5,"['10.1080/0263493032000053208', '10.1007/978-981-13-6693-2_5', 'full/10.1080/09668136.2020.1844867', '10.1038/s41467-020-19493-3', '10.1017/s0020743800021954', None, None, None, '33293507', None, None, None, None, '7723057', None]","[['[[central asian survey'], ['springer singapore'], ['europe-asia studies'], ['nature communications'], ['international journal of middle east studies']]",63,19,0,103,0,4,98,0.21649484536082475,0.06529209621993128,0.3539518900343643,0.01718213058419244,0.0,0.29896907216494845,5,"['www.census.gov', 'stat.gov', 'www.cia.gov', 'minerals.usgs.gov', 'state.gov', '2009-2017.state.gov', 'www.cia.gov', 'whitehouse.gov', 'www.stat.gov', 'www.cia.gov', 'webarchive.loc.gov', '2009-2017.state.gov', 'whitehouse.gov', 'stat.gov', '2009-2017.state.gov', 'www.cia.gov', '2009-2017.state.gov', '2009-2017.state.gov', 'www.stat.gov', 'books.google.com', 'www.nytimes.com', 'www.tax-news.com', 'worldatlas.com', 'www.ogj.com', 'www.taipeitimes.com', 'www.usnews.com', 'astanatimes.com', 'astanatimes.com', 'www.railwaygazette.com', 'books.google.com', 'www.nytimes.com', 'www.bbc.com', 'astanatimes.com', 'webcache.googleusercontent.com', 'books.google.com', 'www.washingtonpost.com', 'www.iihf.com', 'www.economist.com', 'ey.com', 'www.britannica.com', 'www.reuters.com', 'economictimes.indiatimes.com', 'thediplomat.com', 'marginalrevolution.com', 'thediplomat.com', 'tass.com', 'www.france24.com', 'www.raillynews.com', 'www.ebrd.com', 'www.railwaygazette.com', 'bloomberg.com', 'books.google.com', 'www.nytimes.com', 'www.ft.com', 'www.britannica.com', 'gca.satrapia.com', 'www.tasteatlas.com', 'www.usnews.com', 'books.google.com', 'www.britannica.com', 'huffingtonpost.com', 'www.bbc.com', 'www.flightglobal.com', 'encarta.msn.com', 'astanatimes.com', 'finchannel.com', 'www.fitchratings.com', 'www.aljazeera.com', 'forbes.com', 'www.etymonline.com', '2fwww.ft.com', 'www.iran-daily.com', 'www.kazakhembus.com', 'books.google.com', 'www.bricplusnews.com', 'cis-legislation.com', 'www.britannica.com', 'encarta.msn.com', 'www.reuters.com', 'kazakhstanun.com', 'astanatimes.com', 'www.globalpost.com', 'astanatimes.com', 'latino.foxnews.com', 'www.bbc.com', 'www.france24.com', 'www.weatherbase.com', 'astanatimes.com', 'thediplomat.com', 'astanatimes.com', 'www.iran-daily.com', 'astanatimes.com', 'www.theatlantic.com', 'www.forbes.com', 'astanatimes.com', 'www.economist.com', 'homestead.com', 'astanatimes.com', 'www.washingtonpost.com', 'content.time.com', 'www.railjournal.com', 'astanatimes.com', 'www.iht.com', 'www.aa.com', 'www.bbc.com', 'www.bloomberg.com', 'www.reuters.com', 'www.nytimes.com', 'books.google.com', 'thediplomat.com', 'www.business-standard.com', 'www.bloomberg.com', 'astanatimes.com', 'viranatura.com', 'kazakhstan.orexca.com', 'gca.satrapia.com', 'www.sunkarresources.com', 'cannescorporate.com', 'www.bbc.com', 'books.google.com', 'www.economist.com', 'www.studycountry.com', 'www.atlanticcouncil.org', 'treaties.un.org', 'imf.org', 'www.oic-oci.org', 'www.hrw.org', 'pewforum.org', 'world-nuclear.org', 'www.eurasia.undp.org', 'www.hrw.org', 'oecd.org', 'www.americanbar.org', 'www.hrw.org', 'www.hrw.org', 'www3.weforum.org', 'www.pewforum.org', 'www.oecd.org', 'data.worldjusticeproject.org', 'www.pbs.org', 'globalreligiousfutures.org', 'cdi.org', 'www.baselgovernance.org', 'www.forum18.org', 'www.oecd.org', 'www.americanbar.org', 'www.globalreligiousfutures.org', 'www.eurasianet.org', 'www.irinnews.org', 'www.crisisgroup.org', 'asiecentrale.revues.org', 'www.forum18.org', 'un.org', 'pri.org', 'creativecommons.org', 'www.rferl.org', 'monderusse.revues.org', 'freedomhouse.org', 'imf.org', 'data.worldbank.org', 'www.iea.org', 'rsf.org', 'www.americanbar.org', 'www.osce.org', 'rsf.org', 'data.worldbank.org', 'eurasianet.org', 'eiti.org', 'www.doingbusiness.org', 'wto.org', 'whc.unesco.org', 'www.religions-congress.org', 'www.worldbank.org', 'www.heritage.org', 'hdr.undp.org', 'www.wto.org', 'www.unevoc.unesco.org', 'bank.org', 'www.americanbar.org', 'www.collegeatlas.org', 'hrw.org', 'eurasianet.org', 'www.hrw.org', 'www.religions-congress.org', 'whc.unesco.org', ['[[central asian survey'], ['springer singapore'], ['europe-asia studies'], ['nature communications'], ['international journal of middle east studies']]",16642,Require extended confirmed access (no expiry set),245900,11 May 2001,KoyaanisQatsi ,9801,30,2001-05-11,2001-05,2001
227,227,Early Germanic culture,https://en.wikipedia.org/wiki/Early_Germanic_culture,79,1,"['10.16995/trac2007_131_150', None, None]","[['[[theoretical roman archaeology journal', '[[open library of humanities']]",3,0,0,24,0,0,51,0.0379746835443038,0.0,0.3037974683544304,0.012658227848101266,0.0,0.05063291139240506,1,"['books.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.britannica.com', 'www.libertaddigital.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'de.wikipedia.org', 'catalog.hathitrust.org', 'catalog.hathitrust.org', ['[[theoretical roman archaeology journal', '[[open library of humanities']]",62647273,Allow all users (no expiry set),123842,23 December 2019,Krakkos ,111,7,2019-12-23,2019-12,2019
228,228,Dublin,https://en.wikipedia.org/wiki/Dublin,213,3,"['10.2752/175174411x13088262162631', '10.1016/s0140-6736(02)11281-5', '10.5204/mcj.456', None, '12401247', None, None, None, None]","[['food'], ['the lancet'], ['m']]",7,3,0,51,0,2,147,0.03286384976525822,0.014084507042253521,0.23943661971830985,0.014084507042253521,0.0,0.06103286384976526,3,"['www.dccae.gov', 'www.sanjoseca.gov', 'www.liverpool.gov', 'www.irishexperience.com', 'books.google.com', 'www.irishtimes.com', 'www.irishtimes.com', 'www.weather-atlas.com', 'www.irishtimes.com', 'www.irishtimes.com', 'www.irishtimes.com', 'irishtimes.com', 'www.irishtimes.com', 'www.zyen.com', 'www.irishtimes.com', '2fwww.irishtimes.com', 'www.irishtimes.com', 'www.irishtimes.com', 'cricketarchive.com', 'architectural-review.com', 'www.cricketeurope.com', 'www.irishcentral.com', 'books.google.com', 'www.irishtimes.com', '2fwww.irishtimes.com', 'books.google.com', 'www.smh.com', 'irishtimes.com', 'www.irishtimes.com', 'irishtimes.com', 'citymayors.com', 'www.irishtimes.com', 'archiseek.com', 'www.irishtimes.com', 'www.irishtimes.com', 'everything2.com', 'www.irishtimes.com', 'www.nytimes.com', 'issuu.com', 'books.google.com', 'tomtom.com', 'www.irishtimes.com', 'dublinairport.com', 'www.irishtimes.com', 'www.irishtimes.com', 'visitdublin.com', 'www.irishexaminer.com', 'dailyhomelist.com', 'www.citymayors.com', 'books.google.com', 'issuu.com', 'dublinobserver.com', 'www.irishtimes.com', 'www.irishtimes.com', 'www.jstor.org', 'traveldir.org', 'britishcouncil.org', 'britishcouncil.org', 'www.greatirelandrun.org', 'www.jstor.org', 'www.worldcat.org', ['food'], ['the lancet'], ['m']]",8504,Require administrator access (no expiry set),167326,25 September 2001,Eob ,9433,13,2001-09-25,2001-09,2001
229,229,Stockholm,https://en.wikipedia.org/wiki/Stockholm,122,0,[],[],7,1,0,23,0,0,91,0.05737704918032787,0.00819672131147541,0.1885245901639344,0.0,0.0,0.06557377049180328,0,"['www.gov', 'www.tripadvisor.com', 'stockholmtown.com', 'onetomulti.com', 'www.rd.com', 'www.bbc.com', 'www.foreignpolicy.com', 'books.google.com', 'www.visitstockholm.com', 'books.google.com', 'www.businessweek.com', 'www.oyster.com', 'www.nytimes.com', 'www.businessinsider.com', 'www.atptour.com', 'www.citylab.com', 'inhabitat.com', 'articles.chicagotribune.com', 'stockholmnews.com', 'www.stockholmjazz.com', 'www.railjournal.com', 'books.google.com', 'traveler.nationalgeographic.com', 'articles.chicagotribune.com', 'www.stad.org', 'www.norden.org', 'www.mindat.org', 'www.cforic.org', 'sv.climate-data.org', 'commons.wikimedia.org', 'www.stad.org']",26741,Require administrator access (no expiry set),133513,29 August 2001,Pinkunicorn ,5230,13,2001-08-29,2001-08,2001
230,230,Latvia,https://en.wikipedia.org/wiki/Latvia,274,8,"['10.1038/s41467-020-19493-3', '10.1080/00905992.2013.823391', '10.1002/j.1538-165x.2009.tb00657.x', '10.3390/resources7030058', '10.1080/01629778700000141', '10.1080/01629779900000031', '10.1080/01629770100000191', '33293507', None, None, None, None, None, None, '7723057', None, None, None, None, None, None]","[['nature communications'], ['nationalities papers ', '[[cambridge university press'], [' political science quarterly '], ['resources'], ['journal of baltic studies'], ['journal of baltic studies'], ['journal of baltic studies ']]",31,38,0,45,0,2,151,0.11313868613138686,0.1386861313868613,0.16423357664233576,0.029197080291970802,0.0,0.28102189781021897,7,"['webarchive.loc.gov', 'www.csb.gov', 'www.izm.gov', 'data.stat.gov', 'csb.gov', 'www.daba.gov', '2009-2017.state.gov', 'csb.gov', 'data.csb.gov', 'www.tm.gov', 'csb.gov', 'www.mfa.gov', '2009-2017.state.gov', 'www.mfa.gov', 'www.irs.gov', 'www.futureforum2013.gov', 'www.mfa.gov', 'data.csb.gov', 'www.mod.gov', 'www.mk.gov', '2009-2017.state.gov', 'data1.csb.gov', 'data.csb.gov', 'www.csb.gov', 'www.cia.gov', 'www.mfa.gov', 'apps.fas.usda.gov', 'www.csb.gov', 'www.am.gov', 'www.cia.gov', 'www.csb.gov', 'data.csb.gov', '2009-2017.state.gov', 'mod.gov', 'data.csb.gov', 'data.stat.gov', 'www.csb.gov', 'csb.gov', 'www.bbc.com', 'espn.com', 'graphics.eiu.com', 'www.dw.com', 'www.bbc.com', 'www.bayefsky.com', 'www.latimes.com', 'www.lonelyplanet.com', 'www.nytimes.com', 'books.google.com', 'www.history.com', 'www.bloomberg.com', 'www.airbaltic.com', 'onlatvia.com', 'www.defensenews.com', 'bnn-news.com', 'onlatvia.com', 'latviansongfest.com', 'www.nytimes.com', 'www.bbc.com', 'www.washingtonpost.com', 'www.wsj.com', 'flaglog.com', 'www.bbc.com', 'www.baltic-course.com', 'riga-jurmala.com', 'books.google.com', 'www.interkultur.com', 'uefa.com', 'www.baltic-course.com', 'www.lonelyplanet.com', 'healthcare-in-europe.com', 'nhl.com', 'www.reuters.com', 'www.economist.com', 'books.google.com', 'www.balticsworldwide.com', 'findarticles.com', 'www.baltic-course.com', 'www.travelsignposts.com', 'books.google.com', 'lonelyplanet.com', 'books.google.com', 'mongabay.com', 'www.reuters.com', 'www.unhcr.org', 'en.unesco.org', 'stats.oecd.org', 'www.globalsecurity.org', 'www.nordplusonline.org', 'openknowledge.worldbank.org', 'imf.org', 'www.unece.org', 'report2009.amnesty.org', 'www.railbaltica.org', 'www.privacyinternational.org', 'www.lhnet.org', 'www.oecd.org', 'www.nb8businessmobility.org', 'data.footprintnetwork.org', 'www.hrw.org', 'web.worldbank.org', 'www.historyofwar.org', 'www.imc-cim.org', 'www.imf.org', 'www.ndpculture.org', 'www.freedomhouse.org', 'latvianart.org', 'www.gwp.org', 'www.kulturkontaktnord.org', 'hdr.undp.org', 'hdr.undp.org', 'www.europeanfilmacademy.org', 'en.rsf.org', 'web.worldbank.org', 'wayback.archive-it.org', ['nature communications'], ['nationalities papers ', '[[cambridge university press'], [' political science quarterly '], ['resources'], ['journal of baltic studies'], ['journal of baltic studies'], ['journal of baltic studies ']]",17514,Require administrator access (no expiry set),181995,1 March 2001,Josh Grosse ,7375,14,2001-03-01,2001-03,2001
231,231,Nagpur,https://en.wikipedia.org/wiki/Nagpur,356,0,[],[],20,31,0,221,0,0,84,0.056179775280898875,0.08707865168539326,0.6207865168539326,0.0,0.0,0.14325842696629212,0,"['www.nmcnagpur.gov', 'nagpur.gov', 'www.maharashtra.gov', 'www.trai.gov', 'mpsp.maharashtra.gov', 'imdnagpur.gov', 'nagpur.gov', 'mahades.maharashtra.gov', 'census.gov', 'imdpune.gov', 'employmentnews.gov', 'nagpurpolice.gov', 'mp.gov', 'nmcnagpur.gov', 'mpcb.gov', 'mahapolice.gov', 'imdpune.gov', 'www.censusindia.gov', 'cr.indianrailways.gov', 'www.maharashtratourism.gov', 'dcmsme.gov', 'www.nmcnagpur.gov', 'nagpur.gov', 'www.cr.indianrailways.gov', 'allindiaradio.gov', 'imdpune.gov', 'pdf.usaid.gov', 'cr.indianrailways.gov', 'www.cia.gov', 'nagpurpolice.gov', 'www.trai.gov', 'www.nriol.com', 'timesofindia.indiatimes.com', 'zeenews.india.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.thehitavada.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'articles.timesofindia.indiatimes.com', 'www.urbantransportnews.com', 'www.kecrpg.com', 'dwarkapark.com', 'www.infosys.com', 'minexindia.com', 'www.lokmat.com', 'timesofindia.indiatimes.com', 'www.moneycontrol.com', 'www.pixtrans.com', 'www.amuserr.com', 'books.google.com', 'www.suruchiinternational.com', 'www.moneycontrol.com', 'timesofindia.indiatimes.com', 'necoindia.com', 'www.funnfood.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'sanjeevkapoor.com', 'www.bharatcontainers.com', 'nagpur.joiye.com', 'britannica.com', 'www.bhaskar.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'stats.rleague.com', 'www.thehitavada.com', 'timesofindia.indiatimes.com', 'www.highlandparknagpur.com', 'inprotantindia.com', 'articles.timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.thehitavada.com', 'ndtvsports.com', 'books.google.com', 'search.rediff.com', 'www.thehindubusinessline.com', 'books.google.com', 'www.mahamarathon.com', 'books.google.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.kanakresources.com', 'www.mh-31.com', 'www.latestly.com', 'www.hindu.com', 'jain24.com', 'economictimes.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.calderys.com', 'www.holidify.com', 'www.indoramaindia.com', 'mahacid.com', 'www.unitech-power.com', 'timesofindia.indiatimes.com', 'www.firstpost.com', 'www.newindianexpress.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'govtchitrakalamahavidyalayanagpur.com', 'timesofindia.indiatimes.com', 'economictimes.indiatimes.com', 'timesofindia.indiatimes.com', 'www.jointreplacementclinic.com', 'www.thehindu.com', 'economictimes.indiatimes.com', 'timesofindia.indiatimes.com', 'www.cricbuzz.com', 'books.google.com', 'www.thehindu.com', 'www.ocwindia.com', 'timesofindia.indiatimes.com', 'zeenews.india.com', 'www.lokmat.com', 'food.manoramaonline.com', 'timesofindia.indiatimes.com', 'nagpurwater.com', 'thehitavada.com', 'timesofindia.indiatimes.com', '0milemarathon.com', 'indiaelectron.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.deccanherald.com', 'urbantransportnews.com', 'timesofindia.indiatimes.com', 'bombayparsipunchayet.com', 'transrailltd.com', 'www.thehitavada.com', 'financialexpress.com', 'www.business-standard.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.dnaindia.com', 'timesofindia.indiatimes.com', 'nationnext.com', 'timesofindia.indiatimes.com', 'economictimes.indiatimes.com', 'timesofindia.indiatimes.com', 'loksatta.com', 'timesofindia.indiatimes.com', 'fmstations.bharatiyamobile.com', 'zeenews.india.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.livemint.com', 'content-usa.cricinfo.com', 'dnaindia.com', 'www.maidcmumbai.com', 'articles.economictimes.indiatimes.com', 'inprotantindia.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'csridentity.com', 'www.dqweek.com', 'www.ibnlive.com', 'economictimes.indiatimes.com', 'travelspedia.com', 'www.lokmat.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.moneycontrol.com', 'www.poddareshwarrammandir.com', 'timesofindia.indiatimes.com', 'www.amritt.com', 'www.financialexpress.com', 'www.indianexpress.com', 'www.halbadarpan.com', 'timesofindia.indiatimes.com', 'maharashtraweb.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.sanvijay.com', 'timesofindia.indiatimes.com', 'indianexpress.com', 'conferencing.pic.twitter.com', 'www.nagpurorange.com', 'www.business-standard.com', 'articles.economictimes.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'catalign.com', 'timesofindia.indiatimes.com', 'www.deccanchronicle.com', 'www.vccircle.com', 'timesofindia.indiatimes.com', 'buddhistentrepreneurs.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.tribuneindia.com', 'nagpur-hotels.com', 'www.asianage.com', 'www.ibnlive.com', 'thehindu.com', 'timesofindia.indiatimes.com', 'www.mh-31.com', 'www.icc-cricket.com', 'timesofindia.indiatimes.com', 'catalogs.infobanc.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.thehitavada.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.financialexpress.com', 'timesofindia.indiatimes.com', 'www.tribuneindia.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'articles.timesofindia.indiatimes.com', 'hindustantimes.com', 'www.candicoindia.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'food52.com', 'indiansaga.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.hindustantimes.com', 'www.hindu.com', 'jointreplacementclinic.com', 'www.indianexpress.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.firstpost.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.nitnagpur.org', 'www.dmer.org', 'www.nitnagpur.org', 'www.midcindia.org', 'www.unesco.org', 'rchiips.org', 'www.nitnagpur.org', 'www.ddkmumbai.org', 'mls.org', 'download.nos.org', 'rbi.org', 'sangharakshita.org', 'bioanofrontier.org', 'tniusnews.org', 'www.baps.org', 'www.nagpuruniversity.org', 'ijsetr.org', 'indiabiodiversity.org', 'www.india-now.org', 'cbkamptee.org']",460979,Allow all users (no expiry set),178308,8 February 2004,66.69.208.214 ,5703,12,2004-02-08,2004-02,2004
232,232,Albania,https://en.wikipedia.org/wiki/Albania,387,6,"['10.1111/j.1548-1360.2010.01081.x', '10.1038/s41467-020-19493-3', '10.1080/17450101.2012.718939', '10.1657/1938-4246-41.4.455', '10.1093/cje/25.1.1', '10.5209/rev_unis.2011.v26.37824', None, '33293507', None, None, None, None, None, '7723057', None, None, None, None]","[['cultural anthropology '], ['nature communications'], ['mobilities '], ['arctic'], ['cambridge journal of economics '], ['unisci discussion papers ']]",65,47,0,140,0,0,129,0.16795865633074936,0.12144702842377261,0.36175710594315247,0.015503875968992248,0.0,0.3049095607235142,6,"['www.instat.gov', 'ambasadat.gov', 'www.instat.gov', 'state.gov', 'www.instat.gov', 'www.ngdc.noaa.gov', 'www.instat.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', '2009-2017.state.gov', 'www.cia.gov', 'fdi.gov', 'www.instat.gov', 'qbz.gov', 'punetejashtme.gov', 'akzm.gov', 'www.ambasadat.gov', 'mod.gov', 'www.csce.gov', 'www.instat.gov', 'www.instat.gov', 'instat.gov', 'www.qbz.gov', 'www.instat.gov', 'ata.gov', 'shendetesia.gov', '2001-2009.state.gov', 'www.instat.gov', 'shendetesia.gov', 'instat.gov', 'state.gov', 'www.infrastruktura.gov', 'www.export.gov', 'www.moi.gov', 'eia.gov', 'shendetesia.gov', 'www.instat.gov', 'databaza.instat.gov', 'www.cia.gov', 'databaza.instat.gov', 'punetejashtme.gov', 'www.instat.gov', 'www.dsdc.gov', 'www.dfid.gov', 'databaza.instat.gov', 'books.google.com', 'winesofbalkans.com', 'www.balkanchronicle.com', 'books.google.com', 'books.google.com', 'www.bloomberg.com', 'propertywire.com', 'books.google.com', 'books.google.com', 'books.google.com', 'winealbania.com', 'www.britannica.com', 'www.britannica.com', 'books.google.com', 'www.balkaninsight.com', 'books.google.com', 'www.nytimes.com', 'www.ocnal.com', 'balkaneu.com', 'ijbcnet.com', 'www.setimes.com', 'www.britannica.com', 'telegrafi.com', 'referenceworks.brillonline.com', 'books.google.com', 'books.google.com', 'www.tap-ag.com', 'www.panorama.com', 'www.balkanchronicle.com', 'shqiperia.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'shqiptarja.com', 'books.google.com', 'books.google.com', 'books.google.com', 'shekulli.com', 'books.google.com', 'books.google.com', 'shekulli.com', 'shqiptarja.com', 'wingia.com', 'books.google.com', 'books.google.com', 'arkivalajmeve.com', 'books.google.com', 'www.tap-ag.com', 'books.google.com', 'dw.com', 'books.google.com', 'winealbania.com', 'anteacement.com', 'books.google.com', 'books.google.com', 'www.economist.com', 'www.gallup.com', 'novinite.com', 'books.google.com', 'investinmacedonia.com', 'books.google.com', 'albaniainbrief.com', 'www.euronews.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'referenceworks.brillonline.com', 'books.google.com', 'telegrafi.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.ocnal.com', 'dhsprogram.com', 'jacobinmag.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.ethnologue.com', 'www.setimes.com', 'books.google.com', 'nasdaq.com', 'www.ynetnews.com', 'books.google.com', 'books.google.com', 'setimes.com', 'books.google.com', 'books.google.com', 'www.balkaninsight.com', 'www.reuters.com', 'books.google.com', 'books.google.com', 'www.dw.com', 'www.lonelyplanet.com', 'books.google.com', 'www.lonelyplanet.com', 'epicureandculture.com', 'www.worldatlas.com', 'books.google.com', 'macfungi.webs.com', 'books.google.com', 'shekulli.com', 'www.aa.com', 'books.google.com', 'books.google.com', 'tiranatimes.com', 'www.allbusiness.com', 'books.google.com', 'www.travel-gazette.com', 'books.google.com', 'books.google.com', 'forbes.com', 'setimes.com', 'books.google.com', 'books.google.com', 'a2news.com', 'gazeta-shqip.com', 'arkivi.peshkupauje.com', 'shqiptarja.com', 'books.google.com', 'letersia.fajtori.com', 'shqiptarja.com', 'www.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'worldatlas.com', 'theodora.com', 'earthquake-report.com', 'www.newscientist.com', 'www.scribd.com', 'books.google.com', 'www.dw.com', 'www.korrieri.com', 'religion-freedom-report.org', 'rsf.org', 'al.undp.org', 'www.osce.org', 'www.unesco.org', 'www.unocha.org', 'data.worldbank.org', 'biblicalstudies.org', 'osce.org', 'agroweb.org', 'ppnea.org', 'www.imf.org', 'www.undp.org', 'www.imf.org', 'www.gutenberg.org', 'wri-irg.org', 'whc.unesco.org', 'www.ted-adventist.org', 'www.unesco.org', 'www.hydropower.org', 'newsroom.lds.org', 'www.jewishvirtuallibrary.org', 'data.worldbank.org', 'whc.unesco.org', 'osce.org', 'wttc.org', 'ich.unesco.org', 'www.osce.org', 'unece.org', 'invest-in-albania.org', 'ateistet.org', 'www.osce.org', 'faostat.fao.org', 'www.unhcr.org', 'osce.org', 'www.thealbaniancinemaproject.org', 'esc.albaniaenergy.org', 'www.wssinfo.org', 'www.al.undp.org', 'meetingorganizer.copernicus.org', 'freedomhouse.org', 'www.energy-community.org', 'climateknowledgeportal.worldbank.org', 'whc.unesco.org', 'linguistlist.org', 'osce.org', 'wttc.org', 'esc.albaniaenergy.org', 'agroweb.org', 'world.bymap.org', 'www.migrationinformation.org', 'unstats.un.org', 'unece.org', 'hdr.undp.org', 'www.revolutionarydemocracy.org', 'www.imf.org', 'hdi.globaldatalab.org', 'invest-in-albania.org', 'osce.org', 'osce.org', 'wayback.archive-it.org', 'whc.unesco.org', 'mirror.undp.org', 'www.catsg.org', 'www.worlddiplomacy.org', ['cultural anthropology '], ['nature communications'], ['mobilities '], ['arctic'], ['cambridge journal of economics '], ['unisci discussion papers ']]",738,Require administrator access (no expiry set),274933,4 November 2001,H.W. ,16291,5,2001-11-04,2001-11,2001
233,233,Assam,https://en.wikipedia.org/wiki/Assam,275,2,"['10.2307/3517004', '10.2307/603683', None, None, None, None]","[['social scientist'], ['journal of the american oriental society']]",32,19,0,117,0,0,105,0.11636363636363636,0.06909090909090909,0.4254545454545455,0.007272727272727273,0.0,0.19272727272727272,2,"['planningcommission.gov', 'www.assamassembly.gov', 'finance.assam.gov', 'www.censusindia.gov', 'www.eia.gov', 'assamaccord.assam.gov', 'censusindia.gov', 'censusindia.gov', 'karimganj.gov', 'karimganj.gov', 'assamaccord.assam.gov', 'www.censusindia.gov', 'censusindia.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'censusindia.gov', 'online.assam.gov', 'www.censusindia.gov', 'nagaon.gov', 'www.thehindu.com', 'www.pratidintime.com', 'www.reuters.com', 'books.google.com', 'books.google.com', 'assamtribune.com', 'm.economictimes.com', 'indianexpress.com', 'www.thehindu.com', 'hinduonnet.com', 'www.thehindu.com', 'www.telegraphindia.com', 'timesofindia.indiatimes.com', 'indianexpress.com', 'www.telegraphindia.com', 'm.hindustantimes.com', 'books.google.com', 'books.google.com', 'm.timesofindia.com', 'www.assamtribune.com', 'ibnlive.in.com', 'www.sentinelassam.com', 'www.sentinelassam.com', 'www.hindustantimes.com', 'assamco.com', 'www.east-himalaya.com', 'books.google.com', 'www.hindu.com', 'm.ndtv.com', 'm.hindustantimes.com', 'economictimes.indiatimes.com', 'indianexpress.com', 'www.telegraphindia.com', 'www.ethnologue.com', 'www.hindustantimes.com', 'zeenews.india.com', 'm.timesofindia.com', 'www.moneycontrol.com', 'www.indiatvnews.com', 'm.ndtv.com', 'www.arunachaltourism.com', 'silchartoday.com', 'www.indiablooms.com', 'www.assamtribune.com', 'www.sentinelassam.com', 'www.languagesgulper.com', 'm.timesofindia.com', 'www.thehindu.com', 'books.google.com', 'www.ndtv.com', 'www.hindustantimes.com', 'timesofindia.indiatimes.com', 'indianexpress.com', 'books.google.com', 'www.bharatonline.com', 'www.business-standard.com', 'books.google.com', 'www.hindustantimes.com', 'www.hindustantimes.com', 'indianexpress.com', 'www.thehindu.com', 'm.timesofindia.com', 'databank.nedfi.com', 'indianexpress.com', 'books.google.com', 'm.ndtv.com', 'thekararnivang.com', 'm.firstpost.com', 'www.thethumbprintmag.com', 'www.financialexpress.com', 'www.bordowathan.com', 'www.thehindu.com', 'm.economictimes.com', 'www.assamtribune.com', 'timesofindia.indiatimes.com', 'www.business-standard.com', 'm.hindustantimes.com', 'm.hindustantimes.com', 'www.ethnologue.com', 'www.bbc.com', 'thekararnivang.com', 'www.assamtribune.com', 'indiarailinfo.com', 'www.nytimes.com', 'www.newslaundry.com', 'www.assamtribune.com', 'www.hindustantimes.com', 'm.hindustantimes.com', 'm.firstpost.com', 'www.newindianexpress.com', 'investinassam.com', 'www.deccanherald.com', 'www.firstpost.com', 'www.assamtribune.com', 'indiarailinfo.com', 'www.ndtv.com', 'www.assamtribune.com', 'www.news18.com', 'www.thethumbprintmag.com', 'databank.nedfi.com', 'zeenews.india.com', 'www.telegraphindia.com', 'www.thehindu.com', 'm.timesofindia.com', 'www.aljazeera.com', 'www.newindianexpress.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.business-standard.com', 'iloveindia.com', 'books.google.com', 'www.india.com', 'timesofindia.indiatimes.com', 'www.telegraphindia.com', 'www.telegraphindia.com', 'm.timesofindia.com', 'articles.economictimes.indiatimes.com', 'www.assamtourism.org', 'www.dhubrimb.org', 'www.satp.org', 'cdpsindia.org', 'milaap.org', 'bodolanduniversity.org', 'www.envisassam.org', 'faostat.fao.org', 'planassam.org', 'www.alterinter.org', 'satp.org', 'assamgov.org', 'hdi.globaldatalab.org', 'www.downtoearth.org', 'voi.org', 'dibrugarhmunicipality.org', 'www.satp.org', 'www.satp.org', 'milaap.org', 'www.jstor.org', 'goalparamb.org', 'planassam.org', 'satp.org', 'whc.unesco.org', 'www.adb.org', 'www.indiatea.org', 'jorhatmunicipalboard.org', 'www.assamtimes.org', 'en.banglapedia.org', 'www.birdlife.org', 'www.envisassam.org', 'dibrugarhmunicipality.org', ['social scientist'], ['journal of the american oriental society']]",186162,"Require autoconfirmed or confirmed access (18:42, 1 July 2022)",202049,21 February 2003,203.200.38.93 ,8091,24,2003-02-21,2003-02,2003
234,234,Korea,https://en.wikipedia.org/wiki/Korea,224,3,"['10.1007/s10680-005-6851-6', '10.1111/j.1728-4457.2012.00475.x', '10.1177/095624780401600112', None, None, None, None, None, None]","[[' european journal of population '], [' population and development review '], ['environment and urbanization ']]",14,7,0,143,0,0,57,0.0625,0.03125,0.6383928571428571,0.013392857142857142,0.0,0.10714285714285714,3,"['www.cia.gov', 'www.loc.gov', 'www.cia.gov', 'www.loc.gov', 'lcweb2.loc.gov', 'www.loc.gov', '2001-2009.state.gov', 'books.google.com', 'www.japan-guide.com', 'books.google.com', 'english.chosun.com', 'books.google.com', 'books.google.com', 'japan.com', 'books.google.com', 'www.lifeinkorea.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.kimsoft.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', '100.naver.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.everyculture.com', 'books.google.com', 'books.google.com', 'www.everyculture.com', 'msnbc.msn.com', 'www.everyculture.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.oxfordreference.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.japan-guide.com', 'books.google.com', 'books.google.com', 'books.google.com', 'uk.encarta.msn.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.youtube.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.asiasocietymuseum.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thearda.com', 'www.oed.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.atimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'www.aljazeera.com', 'books.google.com', 'books.google.com', 'www.culturecontent.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.newsweek.com', 'books.google.com', 'books.google.com', 'books.google.com', 'news.nationalgeographic.com', 'books.google.com', 'news.naver.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.youtube.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.everyculture.com', 'books.google.com', 'books.google.com', 'www.rightreading.com', 'books.google.com', 'books.google.com', 'news.chosun.com', 'books.google.com', 'www.thoughtco.com', 'books.google.com', 'books.google.com', 'encarta.msn.com', 'books.google.com', 'books.google.com', 'books.google.com', 'articles.latimes.com', 'books.google.com', 'www.oxfordreference.com', 'books.google.com', 'books.google.com', 'encarta.msn.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thoughtco.com', 'www.usnews.com', 'www.bartleby.com', 'books.google.com', 'books.google.com', 'whc.unesco.org', 'whc.unesco.org', 'www.pureinsight.org', 'www.asianinfo.org', 'www.han.org', 'www.metmuseum.org', 'www.nknews.org', 'stats.uis.unesco.org', 'imf.org', 'www.comfort-women.org', 'www.pewforum.org', 'www.metmuseum.org', 'www.oecd.org', 'www.metmuseum.org', [' european journal of population '], [' population and development review '], ['environment and urbanization ']]",16749,Require administrator access (no expiry set),142483,20 July 2001,Andre Engels ,12119,1,2001-07-20,2001-07,2001
235,235,South Korea,https://en.wikipedia.org/wiki/South_Korea,477,6,"['10.1093/acref/9780199568758.001.0001', '10.1038/s41467-020-19493-3', '10.1080/10163270209464030', '10.1017/s1049096510000727', '10.1093/biosci/bix014', None, '33293507', None, None, '28608869', None, '7723057', None, None, '5451287']","[['oxford university press'], ['nature communications'], ['man-ho heo'], ['ps'], ['bioscience']]",55,11,0,224,0,5,176,0.11530398322851153,0.023060796645702306,0.469601677148847,0.012578616352201259,0.0,0.1509433962264151,5,"['www.loc.gov', 'www.cia.gov', 'www.cia.gov', 'www.loc.gov', '2009-2017.state.gov', 'tiq.qld.gov', 'eng.mod.gov', 'www.ustr.gov', 'www.cia.gov', 'www.cia.gov', 'www.ssa.gov', 'books.google.com', 'monitor.icef.com', 'books.google.com', 'www.ameinfo.com', 'www.bbc.com', 'books.google.com', 'www.wsj.com', 'news.chosun.com', 'latimes.com', 'www.nytimes.com', 'www.nytimes.com', 'www.bbc.com', 'www.newsweek.com', 'www.armkor.com', 'www.theatlantic.com', 'books.google.com', 'news.chosun.com', 'www.spacedaily.com', 'www.globalfirepower.com', 'books.google.com', 'www.saveourschools.com', 'www.wingia.com', 'www.upi.com', 'joongangdaily.joins.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.reuters.com', 'fuelcelltoday.com', 'english.chosun.com', 'www.defenseindustrydaily.com', 'books.google.com', 'articles.latimes.com', 'english.chosun.com', 'books.google.com', 'www.newsweek.com', 'books.google.com', 'books.google.com', 'www.straitstimes.com', 'www.thefreelibrary.com', 'fortune.com', 'beyondhallyu.com', 'www.reuters.com', 'books.google.com', 'theconversation.com', 'books.google.com', 'www.supersport.com', 'books.google.com', 'www.reuters.com', 'www.techspot.com', 'news.nationalgeographic.com', 'books.google.com', 'www.atimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'city.udn.com', 'books.google.com', 'www.brecorder.com', 'content.time.com', 'www.nytimes.com', 'books.google.com', 'www.innovationiseverywhere.com', 'www.livescience.com', 'english.chosun.com', 'www.fiercepharma.com', 'english.chosun.com', 'asiatimes.com', 'www.koreaherald.com', 'www.mcgilltribune.com', 'books.google.com', 'nocamels.com', 'www.weareteachers.com', 'books.google.com', 'books.google.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'www.forbes.com', 'english.chosun.com', 'www.usatoday.com', 'books.google.com', 'books.google.com', 'www.voanews.com', 'www.csmonitor.com', 'books.google.com', 'www.koreaherald.com', 'books.google.com', 'books.google.com', 'dsc.discovery.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.formula1.com', 'books.google.com', 'www.nytimes.com', 'theconversation.com', 'english.chosun.com', 'fuelcellseminar.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.apnews.com', 'm.economictimes.com', 'www.washingtonpost.com', 'keepeek.com', 'books.google.com', 'greentechmedia.com', 'keepeek.com', 'books.google.com', 'cnn.com', 'www.economist.com', 'books.google.com', 'joongangdaily.joins.com', 'edition.cnn.com', 'joongangdaily.joins.com', 'books.google.com', 'www.economist.com', 'sthelepress.com', 'www.aljazeera.com', 'www.tradingmarkets.com', 'pt.scribd.com', 'books.google.com', 'english.chosun.com', 'modernkoreanhistory.weebly.com', 'books.google.com', 'www.defencetalk.com', 'uk.reuters.com', 'books.google.com', 'edition.cnn.com', 'koreajoongangdaily.joins.com', 'books.google.com', 'books.google.com', 'joongangdaily.joins.com', 'www.britannica.com', 'content.time.com', 'thediplomat.com', 'books.google.com', 'thediplomat.com', 'www.popsci.com', 'www.thejakartaglobe.com', 'airlineweekly.com', 'graphics.eiu.com', 'blogs.wsj.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.reuters.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.bloomberg.com', 'books.google.com', 'books.google.com', 'thediplomat.com', 'books.google.com', 'www.christianitytoday.com', 'books.google.com', 'books.google.com', 'books.google.com', 'kushibo.blogspot.com', 'books.google.com', 'books.google.com', 'www.nationmaster.com', 'dynamic-korea.com', 'books.google.com', 'www.businessinsider.com', 'books.google.com', 'deadline.com', 'books.google.com', 'qz.com', 'article.joins.com', 'alhockey.com', 'www.youtube.com', 'www.koreanair.com', 'books.google.com', 'news.xinhuanet.com', 'www.economist.com', 'www.nytimes.com', 'www.bloomberg.com', 'www.nytimes.com', 'books.google.com', 'www.scmp.com', 'www.newsweek.com', 'cnn.com', 'terms.naver.com', 'books.google.com', 'www.google.com', 'news.naver.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'www.theverge.com', 'latimesblogs.latimes.com', 'english.chosun.com', 'www.nytimes.com', 'atimes.com', 'www.upi.com', 'books.google.com', 'books.google.com', 'www.amazon.com', 'www.nationalgeographic.com', 'www.reuters.com', 'nasaspaceflight.com', 'www.nytimes.com', 'books.google.com', 'www.nytimes.com', 'theconversation.com', 'www.reuters.com', 'books.google.com', 'www.nationmultimedia.com', 'www.buddhismtoday.com', 'worldpoliticsreview.com', 'books.google.com', 'www.dokdo-takeshima.com', 'books.google.com', 'www.universityworldnews.com', 'www.forbes.com', 'books.google.com', 'joongangdaily.joins.com', 'www.asiafoundation.org', 'www.oecd.org', 'www.comfort-women.org', 'www.jpri.org', 'npr.org', 'www.oecd.org', 'data.worldbank.org', 'www.imf.org', 'www.umdcipe.org', 'siteresources.worldbank.org', 'imf.org', 'www.asianinfo.org', 'www.imf.org', 'www.christenseninstitute.org', 'gpseducation.oecd.org', 'www3.weforum.org', 'www.oecdbetterlifeindex.org', 'gpseducation.oecd.org', 'data.oecd.org', 'daccess-dds-ny.un.org', 'globalsecurity.org', 'worldbank.org', 'park.org', 'rsf.org', 'www.oecd.org', 'koreandrama.org', 'data.worldbank.org', 'www.globalsecurity.org', 'www.asianinfo.org', 'www.npr.org', 'www.globalsecurity.org', 'globalsecurity.org', 'www.imf.org', 'www.world-nuclear-news.org', 'apexart.org', 'hdr.undp.org', 'www.asianinfo.org', 'transparency.org', 'www.armscontrol.org', 'www.metmuseum.org', 'www.wtf.org', 'stats.oecd.org', 'nobelprize.org', 'bio2008.org', 'www.pri.org', 'www.oecdbetterlifeindex.org', 'www.iter.org', 'www.asianinfo.org', 'gpseducation.oecd.org', 'ich.unesco.org', 'whc.unesco.org', 'www.pri.org', 'globalsecurity.org', 'www.welfareasia.org', 'seoul.triathlon.org', ['oxford university press'], ['nature communications'], ['man-ho heo'], ['ps'], ['bioscience']]",27019,Require administrator access (no expiry set),285643,8 July 2001,TimShell ,19996,27,2001-07-08,2001-07,2001
236,236,Munich,https://en.wikipedia.org/wiki/Munich,138,2,"['10.1038/d41586-018-07208-0', '10.1016/j.tmp.2017.09.003', '30382228', None, None, None]","[['nature '], ['tourism management perspectives ']]",1,2,0,28,0,0,105,0.007246376811594203,0.014492753623188406,0.2028985507246377,0.014492753623188406,0.0,0.036231884057971016,2,"['www.edinburgh.gov', 'www.edinburgh.gov', 'oktoberfestbeerfestivals.com', 'www.panaceapublishinginternational.com', 'munichfound.com', 'books.google.com', 'www.viamichelin.com', 'munichfound.com', 'www.weatherbase.com', 'mobilityexchange.mercer.com', 'www.com', 'riverbreak.com', 'paulaner-nockherberg.com', 'traveler.nationalgeographic.com', 'www.spottedbylocals.com', 'www.youtube.com', 'verona.com', 'www.mercer.com', 'www.inside-munich.com', 'www.destination-munich.com', 'www.inside-munich.com', '2fgo.gale.com', 'paulaner-nockherberg.com', 'money.cnn.com', 'moovitapp.com', 'www.toytowngermany.com', 'www.forbes.com', 'gamesbids.com', 'moovitapp.com', 'www.mercerhr.com', 'www.openrailwaymap.org', ['nature '], ['tourism management perspectives ']]",19058,Allow all users (no expiry set),175022,19 October 2001,Paul Drye ,6634,6,2001-10-19,2001-10,2001
237,237,Gastronationalism,https://en.wikipedia.org/wiki/Gastronationalism,27,5,"['10.1007/s10460-006-9003-7', '10.23943/princeton/9780691154930.003.0003', '10.1017/nps.2019.104', '10.1177/0003122410372226', '10.1002/9780470670590.wbeog226', None, None, None, None, None, None, None, None, None, None]","[['[[agriculture and human values'], ['[[princeton university press'], ['nationalities papers', '[[cambridge university press'], ['[[american sociological review'], ['john wiley ']]",4,0,0,10,0,0,8,0.14814814814814814,0.0,0.37037037037037035,0.18518518518518517,0.0,0.3333333333333333,5,"['www.thestar.com', 'aljazeera.com', 'www.nbcnews.com', 'chopinandmysaucepan.com', 'www.bbc.com', 'www.sbs.com', 'www.scmp.com', 'books.google.com', 'www.borgenmagazine.com', 'asiancorrespondent.com', 'www.worldcat.org', 'www.npr.org', 'www.worldcat.org', 'www.worldcat.org', ['[[agriculture and human values'], ['[[princeton university press'], ['nationalities papers', '[[cambridge university press'], ['[[american sociological review'], ['john wiley ']]",68554701,Allow all users (no expiry set),24844,24 August 2021,Valereee ,83,0,2021-08-24,2021-08,2021
238,238,Cyprus,https://en.wikipedia.org/wiki/Cyprus,284,8,"['10.21773/boun.25.2.6', '10.5194/hess-11-1633-2007', '10.1038/s41467-020-19493-3', '10.1080/10408398209527361', '10.5325/jeasmedarcherstu.3.2.0128', '10.1093/biosci/bix014', '10.1080/0275720032000136642', '10.1111/j.1529-8817.2005.00224.x', None, None, '33293507', '6337782', None, '28608869', None, '16626331', None, None, '7723057', None, None, '5451287', None, None]","[['bogazici journal '], ['hydrol. earth syst. sci. '], ['nature communications '], ['crc critical reviews in food science and nutrition '], ['journal of eastern mediterranean archaeology '], ['bioscience '], ['history and anthropology '], [' annals of human genetics']]",26,27,0,109,0,2,112,0.09154929577464789,0.09507042253521127,0.38380281690140844,0.028169014084507043,0.0,0.2147887323943662,8,"['2009-2017.state.gov', 'www.nam.gov', 'www.moa.gov', 'www.cia.gov', 'www.cia.gov', 'lcweb2.loc.gov', 'www.mof.gov', 'www.cyprus.gov', 'cia.gov', 'cyprus.gov', 'www.cyprus.gov', 'www.loc.gov', 'www.moa.gov', 'www.cyprus.gov', 'www.cia.gov', 'www.moi.gov', 'www.mfa.gov', 'www.metoffice.gov', 'www.moa.gov', 'mcw.gov', 'lcweb2.loc.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.cystat.gov', 'www.presidency.gov', 'www.presidency.gov', 'books.google.com', 'books.google.com', 'www.hurriyetdailynews.com', 'books.google.com', 'books.google.com', 'books.google.com', 'worldpopulationreview.com', 'books.google.com', 'apropertyincyprus.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.reuters.com', 'books.google.com', 'books.google.com', 'www.filmbirth.com', 'books.google.com', 'jacobinmag.com', 'books.google.com', 'cyprus-mail.com', 'www.reuters.com', 'www.philatelism.com', 'www.hurriyetdailynews.com', 'books.google.com', 'famagusta-gazette.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.cyprusbybus.com', 'www.artnet.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'books.google.com', 'geosite.jankrogh.com', 'urban-keys.com', 'books.google.com', 'www.middle-east-confidential.com', 'books.google.com', 'books.google.com', 'greekreporter.com', 'www.worldatlas.com', 'urban-keys.com', 'www.weather2travel.com', 'www.stratfor.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.time.com', 'www.worldatlas.com', 'books.google.com', 'www.philatelism.com', 'books.google.com', 'edition.cnn.com', 'books.google.com', 'www.frieze.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'cyprusbadminton.com', 'www.iht.com', 'books.google.com', 'palaeolexicon.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.aljazeera.com', 'www.apnewsarchive.com', 'www.euroasia-interconnector.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.reuters.com', 'books.google.com', 'travel.nationalgeographic.com', 'www.cyprus-mail.com', 'books.google.com', 'hurarsiv.hurriyet.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.ekathimerini.com', 'www.cyprus-mail.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.iht.com', 'www.worldatlas.com', 'books.google.com', 'www.aljazeera.com', 'books.google.com', 'www.philatelism.com', 'books.google.com', 'books.google.com', 'www.imf.org', 'www.asor.org', 'www.globalreligiousfutures.org', 'www.freedomhouse.org', 'childinfo.org', 'www.imf.org', 'diko.org', 'data.worldbank.org', 'www.imf.org', 'www.crisisgroup.org', 'freedomhouse.org', 'nufussayimi.devplan.org', 'www.imf.org', 'www.cyprusun.org', 'www.prio.org', 'www.globalreligiousfutures.org', 'unstats.un.org', 'hdr.undp.org', 'hdr.undp.org', 'index.rsf.org', 'www.un.org', 'esa.un.org', 'ohchr.org', 'wayback.archive-it.org', 'www.crisisgroup.org', 'data.worldbank.org', ['bogazici journal '], ['hydrol. earth syst. sci. '], ['nature communications '], ['crc critical reviews in food science and nutrition '], ['journal of eastern mediterranean archaeology '], ['bioscience '], ['history and anthropology '], [' annals of human genetics']]",5593,Require administrator access (no expiry set),207947,2 November 2001,193.133.134.xxx ,13483,11,2001-11-02,2001-11,2001
239,239,Bengali Hindus,https://en.wikipedia.org/wiki/Bengali_Hindus,155,5,"['10.1525/gfc.2010.10.3.58', '10.1163/15685270252772759', '10.2307/3516391', '10.1017/s0041977x00112418', None, '10.1163/2589742x-00601003', None, None, None, None, None, None, None, None, None, None, None, None]","[['gastronomica'], ['numen'], ['social scientist'], ['bulletin of the school of oriental and african studies'], ['proceedings of the indian history congress'], ['journal of religion and demography']]",9,2,0,69,0,0,69,0.05806451612903226,0.012903225806451613,0.44516129032258067,0.03225806451612903,0.0,0.1032258064516129,6,"['www.censusindia.gov', 'www.censusindia.gov', 'encyclopedia2.thefreedictionary.com', 'timesofindia.indiatimes.com', 'books.google.com', 'timesofindia.indiatimes.com', 'indianewsrepublic.com', 'frontline.thehindu.com', 'www.dhakatribune.com', 'books.google.com', 'www.dailypioneer.com', 'books.google.com', 'economictimes.indiatimes.com', 'www.nationalheraldindia.com', 'www.magzter.com', 'articles.timesofindia.indiatimes.com', 'archive.indianexpress.com', 'www.trtworld.com', 'www.hindustantimes.com', 'economictimes.indiatimes.com', 'www.telegraphindia.com', 'www.thehindu.com', 'www.aljazeera.com', 'www.timesnownews.com', 'www.odiakitchen.com', 'articles.timesofindia.indiatimes.com', 'www.asianage.com', 'www.aljazeera.com', 'books.google.com', 'www.outlookindia.com', 'indianonlinepages.com', 'timesofindia.indiatimes.com', 'theculturetrip.com', 'www.news18.com', 'books.google.com', 'garamchai.com', 'timesofindia.indiatimes.com', 'gradworks.umi.com', 'www.thehindu.com', 'discovermagazine.com', 'www.oxfordbibliographies.com', 'www.telegraphindia.com', 'www.anandabazar.com', 'www.bbc.com', 'www.firstpost.com', 'www.thestatesman.com', 'www.nytimes.com', 'books.google.com', 'www.expressindia.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'theculturetrip.com', 'indianexpress.com', 'www.radianceweekly.com', 'www.globalfront.com', 'books.google.com', 'www.populationu.com', 'www.exploreandaman.com', 'www.outlookindia.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.outlookindia.com', 'magazine.outlookindia.com', 'www.hindustantimes.com', 'books.google.com', 'outlookindia.com', 'books.google.com', 'www.thecanadianencyclopedia.com', 'www.outlookindia.com', 'www.telegraphindia.com', 'www.kaladanpress.org', 'www.banglastories.org', 'www.londonkalibari.org', 'hdr.undp.org', 'www.indopedia.org', 'www.rabindra-rachanabali.nltr.org', 'www.migrationinformation.org', 'www.jstor.org', 'puja.org', ['gastronomica'], ['numen'], ['social scientist'], ['bulletin of the school of oriental and african studies'], ['proceedings of the indian history congress'], ['journal of religion and demography']]",28003496,Allow all users (no expiry set),89984,11 July 2010,BengaliHindu ,1618,8,2010-07-11,2010-07,2010
240,240,Gold,https://en.wikipedia.org/wiki/Gold,209,40,"['10.1088/2041-8205/774/2/l23', '10.1006/biol.1997.0123', '10.1111/j.1365-2044.1986.tb12920.x', '10.1021/cr980431o', '10.1016/0375-6742(88)90051-9', '10.2478/s13531-011-0052-3', '10.1007/s10787-007-0021-x', '10.1002/9783527633104.ch7', '10.1211/jpp.60.8.0005', '10.1515/9783110470734-013', '10.1016/0019-2791(71)90496-4', '10.1086/190111', '10.1103/physrevb.6.4370', '10.1038/nature10399', '10.1016/j.chemphys.2004.09.023', '10.1080/00207450212018', '10.1034/j.1600-0536.2001.440107-22.x', '10.1039/b708844m', '10.1103/physrevb.77.155401', '10.1126/science.290.5489.117', '10.1007/bf01505547', '10.1038/500535a', '10.1016/j.solidstatesciences.2005.06.015', '10.1081/clt-100108516', '10.2903/j.efsa.2016.4362', '10.1038/s41467-017-00821-z', '10.1080/14686996.2019.1585145', '10.1111/j.1945-5100.1997.tb01242.x', '10.1103/physrev.60.473', '10.1177/28.1.6153194', '10.1002/ange.19270401103', '10.1002/anie.200600274', '10.1016/0012-821x(90)90060-b', '10.1016/0040-1951(90)90089-q', '10.1038/376238a0', '10.1016/j.jclepro.2012.01.042', '10.1103/physrevc.23.1044', '10.1086/203868', '10.1002/1521-3749(200109)627:9<2112::aid-zaac2112>3.0.co;2-2', None, '9637749', '3022615', '11749494', None, None, '18523733', None, '18644191', '29394026', '4110101', None, None, '21901010', None, '12152404', '11156030', '18762832', None, '11021792', None, '23985867', None, '11778673', None, '29018198', '30956731', None, None, '6153194', None, '16639770', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, '5634996', '6442207', None, None, None, None, None, None, None, None, None, None, None, None]","[['the astrophysical journal letters '], ['biologicals '], ['anaesthesia '], ['chemical reviews '], ['journal of geochemical exploration '], ['central european journal of engineering '], ['inflammopharmacology '], ['wiley-vch verlag gmbh '], ['journal of pharmacy and pharmacology '], ['metal ions in life sciences '], ['immunochemistry'], ['the astrophysical journal supplement series '], ['physical review b '], ['nature '], ['chemical physics '], ['the international journal of neuroscience '], ['contact dermatitis '], ['chemical society reviews '], ['physical review b'], ['science '], ['die naturwissenschaften '], ['[[nature '], ['solid state sciences '], ['clinical toxicology '], ['efsa journal '], ['nature communications '], ['sci. technol. adv. mater. '], ['meteoritics '], ['[[physical review'], ['journal of histochemistry and cytochemistry '], ['zeitschrift für angewandte chemie'], ['angewandte chemie international edition '], ['earth and planetary science letters '], ['tectonophysics '], ['nature '], ['journal of cleaner production '], ['[[physical review c'], ['current anthropology '], ['journal of inorganic and general chemistry ']]",16,6,0,94,0,1,52,0.07655502392344497,0.028708133971291867,0.44976076555023925,0.19138755980861244,0.0,0.2966507177033493,39,"['minerals.usgs.gov', 'www.food.gov', 'www.nzpam.gov', 'library.lanl.gov', 'www.nndc.bnl.gov', 'epubs.nsla.nv.gov', 'deseretnews.com', 'books.google.com', 'www.oxfordislamicstudies.com', 'superiormining.com', 'books.google.com', 'www.epicurious.com', 'books.google.com', 'americansilvereagletoday.com', 'www.delafee.com', 'www.kodak.com', 'www.espi-metals.com', 'www.utilisegold.com', 'www.bbc.com', 'www.sciencedaily.com', 'www.marketwatch.com', 'www.wsj.com', 'ausbullion.blogspot.com', 'books.google.com', 'www.smithsonianmag.com', 'www.nytimes.com', 'www.nytimes.com', 'kitco.com', 'books.google.com', 'www.sierranevadavirtualmuseum.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'www.kitco.com', 'books.google.com', 'books.google.com', 'www.highbeam.com', 'books.google.com', 'books.google.com', 'scientificamerican.com', 'apnews.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'www.technology.matthey.com', 'books.google.com', 'books.google.com', 'news.yahoo.com', 'books.google.com', 'www.oxfordislamicstudies.com', 'books.google.com', 'www.marketwatch.com', 'portaracqg.com', 'www.bloomberg.com', 'www.nytimes.com', 'books.google.com', 'www.mining-technology.com', 'chemistry.about.com', 'books.google.com', 'books.google.com', 'oilprice.com', 'www.gold-eagle.com', 'books.google.com', 'scribd.com', 'www.ameinfo.com', 'www.wsj.com', 'news.coinupdate.com', 'www.kitco.com', 'www.cnbc.com', 'medium.com', 'arizonagoldprospectors.com', 'afrinik.com', 'www.popsci.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.cosmosmagazine.com', 'books.google.com', 'www.reuters.com', 'www.investopedia.com', 'www.tanaka-precious.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'www.usfunds.com', 'www.reuters.com', 'www.efgbank.com', 'www.smithsonianmag.com', 'www.forexyard.com', 'www.techradar.com', 'geology.com', 'books.google.com', 'books.google.com', 'ameinfo.com', 'bullionvault.com', 'goldsilver.com', 'www.ligo.org', 'gold.org', 'www.iso.org', 'gold.org', 'www.worstpolluted.org', 'www.goldbulletin.org', 'www.gold.org', 'lbma.org', 'www.nchistoricsites.org', 'www.sciencemag.org', 'www.iisd.org', 'www.unido.org', 'www.gold.org', 'www.webexhibits.org', 'www.usdebtclock.org', 'www.georgiamagazine.org', ['the astrophysical journal letters '], ['biologicals '], ['anaesthesia '], ['chemical reviews '], ['journal of geochemical exploration '], ['central european journal of engineering '], ['inflammopharmacology '], ['wiley-vch verlag gmbh '], ['journal of pharmacy and pharmacology '], ['metal ions in life sciences '], ['immunochemistry'], ['the astrophysical journal supplement series '], ['physical review b '], ['nature '], ['chemical physics '], ['the international journal of neuroscience '], ['contact dermatitis '], ['chemical society reviews '], ['physical review b'], ['science '], ['die naturwissenschaften '], ['[[nature '], ['solid state sciences '], ['clinical toxicology '], ['efsa journal '], ['nature communications '], ['sci. technol. adv. mater. '], ['meteoritics '], ['[[physical review'], ['journal of histochemistry and cytochemistry '], ['zeitschrift für angewandte chemie'], ['angewandte chemie international edition '], ['earth and planetary science letters '], ['tectonophysics '], ['nature '], ['journal of cleaner production '], ['[[physical review c'], ['current anthropology '], ['journal of inorganic and general chemistry ']]",12240,Require administrator access (no expiry set),136114,10 August 2001,Drj ,6932,9,2001-08-10,2001-08,2001
241,241,Culture of Georgia (country),https://en.wikipedia.org/wiki/Culture_of_Georgia_(country),9,0,[],[],0,2,0,0,0,0,7,0.0,0.2222222222222222,0.0,0.0,0.0,0.2222222222222222,0,"['art.gov', 'www.art.gov']",341997,Allow all users (no expiry set),21231,16 October 2003,Lisiate ,503,1,2003-10-16,2003-10,2003
242,242,Cuba,https://en.wikipedia.org/wiki/Cuba,438,24,"['10.2307/20047491', '10.1016/j.eeh.2020.101376', '10.1093/biosci/bix014', '10.1353/jod.0.0051', '10.1111/j.1467-7709.1994.tb00611.x', '10.1177/0169796x19826731', '10.1503/cmaj.1080068', '10.18475/cjos.v43i1.a9', '10.1215/9780822392859', '10.2307/165789', '10.1017/s0022216x0133626x', '10.1017/s0043887120000106', '10.1136/bmj.333.7566.464', '10.1017/s0022216x00012670', '10.1038/s41467-020-19493-3', '10.1080/13683500.2018.1446920', '10.1353/hrq.2007.0033', '10.2307/422443', '10.1080/13510347.2019.1629420', '10.1371/journal.pgen.1004488', '10.1017/s0022216x96004646', '10.1111/laps.12017', '10.1007/s10668-012-9338-8', None, None, '28608869', None, None, None, '18663207', None, None, None, None, None, '16946334', None, '33293507', None, None, None, None, '25058410', None, None, None, None, None, '5451287', None, None, None, '2474886', None, None, None, None, None, '1557950', None, '7723057', None, None, None, None, '4109857', None, None, None]","[[' [[foreign affairs'], ['explorations in economic history'], ['bioscience'], [' journal of democracy '], ['[[society for historians of american foreign relations'], ['journal of developing societies'], ['cmaj '], ['[[caribbean journal of science', 'college of arts and sciences'], ['[[duke university press'], [' [[university of miami'], [' [[journal of latin american studies'], ['world politics'], [' [[bmj'], [' [[journal of latin american studies'], ['nature communications'], ['current issues in tourism'], [' [[human rights quarterly'], ['comparative politics'], ['democratization'], ['plos genetics '], [' journal of latin american studies '], ['latin american politics and society'], ['environment']]",67,18,0,179,0,7,144,0.15296803652968036,0.0410958904109589,0.408675799086758,0.0547945205479452,0.0,0.24885844748858446,23,"['2009-2017.state.gov', 'www.census.gov', 'minerals.usgs.gov', 'www.loc.gov', 'cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'cia.gov', 'www.cia.gov', 'www.fas.usda.gov', 'minerals.usgs.gov', 'www.america.gov', '1997-2001.state.gov', 'www.cia.gov', 'www.america.gov', '2009-2017.state.gov', 'www.goodreads.com', 'www.com', 'iworldnewsservice.com', 'www.reason.com', 'books.google.com', 'www.economist.com', 'www.economist.com', 'books.google.com', 'books.google.com', 'college.cengage.com', 'www.ethnologue.com', 'books.google.com', 'www.nbcnews.com', 'www.miamiherald.com', 'www.afp.com', 'time.com', 'www.cnn.com', 'wsj.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'www.technologyreview.com', 'www.nytimes.com', 'www.poemhunter.com', 'www.nytimes.com', 'www.aljazeera.com', 'economist.com', 'eiu.com', 'www.usatoday.com', 'history.com', 'www.britannica.com', 'moroccotimes.com', 'www.nytimes.com', 'www.latimes.com', 'aljazeera.com', 'themilitant.com', 'www.reference.com', 'whatcuba.com', 'books.google.com', 'www.aljazeera.com', 'www.nytimes.com', 'news.xinhuanet.com', 'www.cnn.com', 'books.google.com', 'www.miamiherald.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'www.nytimes.com', 'www.thecubanhistory.com', 'historytoday.com', 'books.google.com', 'www.usatoday.com', 'abcnews.go.com', 'books.google.com', 'latinostories.com', 'www.usatoday.com', 'www.ethnologue.com', 'books.google.com', 'www.reuters.com', 'edition.cnn.com', 'www.nytimes.com', 'sonentero.blogspot.com', 'www.miamiherald.com', 'www.msn.com', 'www.nationalgeographic.com', 'abcnews.go.com', 'www.bloomberg.com', 'books.google.com', 'books.google.com', 'longitudebooks.com', 'books.google.com', 'www.nytimes.com', 'www.nytimes.com', 'beta.theglobeandmail.com', 'www.politifact.com', 'www.miamiherald.com', 'www.time.com', 'books.google.com', 'fresnoalliance.com', 'www.premierboxingchampions.com', 'aljazeera.com', 'books.google.com', 'semanarioaqui.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.mercatrade.com', 'www.nytimes.com', 'www.washingtonpost.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'about.com', 'books.google.com', 'books.google.com', 'worldpopulationreview.com', 'www.washingtonpost.com', 'www.theatlantic.com', 'books.google.com', 'newspapers.com', 'nationalpost.com', 'www.spanamwar.com', 'www.economist.com', 'aljazeera.com', 'www.reuters.com', 'sports.yahoo.com', 'www.bbc.com', 'books.google.com', 'www.washingtonpost.com', 'www.britannica.com', 'www.washingtonpost.com', 'books.google.com', 'www.nbcnews.com', 'www.efe.com', 'books.google.com', 'www.thepeninsulaqatar.com', 'blog.fonoma.com', 'books.google.com', 'www.bbc.com', 'amp.france24.com', 'books.google.com', 'www.huffingtonpost.com', 'books.google.com', 'books.google.com', 'www.forbes.com', 'voanews.com', 'en.mercopress.com', 'www.reuters.com', 'www.reuters.com', 'books.google.com', 'books.google.com', 'www.ibtimes.com', 'books.google.com', 'datareportal.com', 'www.usatoday.com', 'books.google.com', 'www.sipiapa.com', 'www.nytimes.com', 'whatlatinamerica.com', 'www.arrowsmithpress.com', 'www.nytimes.com', 'books.google.com', 'www.reason.com', 'books.google.com', 'www.cnn.com', 'books.google.com', 'www.nytimes.com', 'popcrush.com', 'warfarehistorynetwork.com', 'www.redorbit.com', 'www.usatoday.com', 'noticias24.com', 'piie.com', 'www.bbc.com', 'www.nbcnews.com', 'www.efe.com', 'www.suenacubano.com', 'books.google.com', 'www.nbcnews.com', 'go.gale.com', 'books.google.com', 'www.afp.com', 'www.rbth.com', 'books.google.com', 'books.google.com', 'www.smithsonianmag.com', 'www.usatoday.com', 'historyofcuba.com', 'books.google.com', 'news.xinhuanet.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.dw.com', 'siteresources.worldbank.org', 'www.pbs.org', 'news.bahai.org', 'www.ascecuba.org', 'dollarsandsense.org', 'arabia.reporters-sans-frontieres.org', 'www.cubacenter.org', 'www.un.org', 'www.latinamericanstudies.org', 'www.hrw.org', 'mdgs.un.org', 'jfklibrary.org', 'www.pewforum.org', 'olympic.org', 'www.constitutionnet.org', 'oxfamamerica.org', 'cfr.org', 'hdr.undp.org', 'index.rsf.org', 'freedomhouse.org', 'www.constitutionnet.org', 'www.cubagenweb.org', 'www.hrw.org', 'news.un.org', 'www.ascecuba.org', 'esa.un.org', 'www.rsf.org', 'www.ascecuba.org', 'openlibrary.org', 'www.jstor.org', 'museodelaresistencia.org', 'www.amnesty.org', 'www.ascecuba.org', 'www.ascecuba.org', 'globalvoicesonline.org', 'www.pbs.org', 'www.todocuba.org', 'www.wola.org', 'millercenter.org', 'alfredcarrada.org', 'www.sipri.org', 'legacy.intracen.org', 'www.ascecuba.org', 'globalsecurity.org', 'www.pbs.org', 'data.worldbank.org', 'www.rsf.org', 'www.hrw.org', 'cubagenweb.org', 'www.un.org', 'www.constituteproject.org', 'www.cidh.org', 'www.refworld.org', 'havanatimes.org', 'rsf.org', 'unstats.un.org', 'www.pbs.org', 'www.guttmacher.org', 'www.rand.org', 'cpj.org', 'www.jstor.org', 'cpj.org', 'www.hrw.org', 'dollarsandsense.org', 'treaties.un.org', 'www.ascecuba.org', 'natcath.org', [' [[foreign affairs'], ['explorations in economic history'], ['bioscience'], [' journal of democracy '], ['[[society for historians of american foreign relations'], ['journal of developing societies'], ['cmaj '], ['[[caribbean journal of science', 'college of arts and sciences'], ['[[duke university press'], [' [[university of miami'], [' [[journal of latin american studies'], ['world politics'], [' [[bmj'], [' [[journal of latin american studies'], ['nature communications'], ['current issues in tourism'], [' [[human rights quarterly'], ['comparative politics'], ['democratization'], ['plos genetics '], [' journal of latin american studies '], ['latin american politics and society'], ['environment']]",5042481,Require administrator access (no expiry set),229702,3 September 2001,Koyaanis Qatsi ,14051,13,2001-09-03,2001-09,2001
243,243,Egyptian cheese,https://en.wikipedia.org/wiki/Egyptian_cheese,23,1,"['10.1128/aem.01667-06', '17189434', '1828670']",[['appl environ microbiol ']],0,0,0,17,0,0,5,0.0,0.0,0.7391304347826086,0.043478260869565216,0.0,0.043478260869565216,1,"['books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'cheese.com', 'books.google.com', ['appl environ microbiol ']]",39109874,Allow all users (no expiry set),16577,14 April 2013,Aymatth2 ,109,0,2013-04-14,2013-04,2013
244,244,Kashmiris,https://en.wikipedia.org/wiki/Kashmiris,16,0,[],[],0,2,0,11,0,0,3,0.0,0.125,0.6875,0.0,0.0,0.125,0,"['www.censusindia.gov', '(.gov', 'tribune.com', 'www.museindia.com', 'books.google.com', 'dawn.com', 'www.britannica.com', 'books.google.com', 'thaindian.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com']",3930749,Allow all users (no expiry set),28993,2 February 2006,Gnikhil ,3095,3,2006-02-02,2006-02,2006
245,245,Ottoman Empire,https://en.wikipedia.org/wiki/Ottoman_Empire,283,21,"['10.1017/s0041977x00149006', '10.1080/01419870701491937', '10.1080/00905990500504871', '10.2143/turc.30.0.2004296', '10.2307/596868', '10.2307/2212668', '10.1353/jwh.2014.0005', '10.1080/14623520801950820', '10.1017/s0007087403005302', '10.1080/15456870.2015.1090439', '10.1080/00263200701422600', '10.1111/0020-8833.00053', '10.1017/s0020743800027276', '10.1086/694391', '10.1177/002182860503600401', '10.4000/monderusse.39', '10.4321/s1130-14732006000200012', '10.1080/00263207908700415', '10.2478/udi-2018-0006', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, '16721484', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None]","[['bulletin of the school of oriental and african studies'], ['ethnic and racial studies '], ['[[nationalities papers'], ['turcica ', 'éditions klincksieck '], ['journal of the american oriental society '], ['the american journal of international law '], ['journal of world history '], ['journal of genocide research '], ['the british journal for the history of science ', '[[cambridge university press'], ['atlantic journal of communication '], ['middle eastern studies '], ['[[international studies quarterly'], ['international journal of middle east studies '], ['the journal of modern history '], ['journal for the history of astronomy ', 'science history publications ltd. '], ['cahiers du monde russe '], ['neurocirugía '], ['middle eastern studies '], ['urban development issues ']]",10,2,0,82,0,1,168,0.0353356890459364,0.007067137809187279,0.28975265017667845,0.07420494699646643,0.0,0.1166077738515901,19,"['www.kultur.gov', 'www.mfa.gov', 'books.google.com', 'warfare.atwebpages.com', 'cache-media.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.howtotalkaboutarthistory.com', 'books.google.com', 'www.twareekh.com', 'www.saudiaramcoworld.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.google.com', 'books.google.com', 'books.google.com', 'global.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'sursockhouse.com', 'www.britannica.com', 'www.oxfordreference.com', 'books.google.com', 'www.emaanlibrary.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'history.com', 'books.google.com', 'books.google.com', 'www.allaboutturkey.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'www.google.com', 'books.google.com', 'history.com', 'www.oxfordislamicstudies.com', 'books.google.com', 'books.google.com', 'www.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.turkeyswar.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'www.google.com', 'books.google.com', 'www.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'global.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.jstor.org', 'www.nationalgeographic.org', 'www.nationalgeographic.org', 'iranicaonline.org', 'faith-matters.org', 'nationalinterest.org', 'globaled.org', 'www.njegos.org', 'historycooperative.org', 'wayback.archive-it.org', ['bulletin of the school of oriental and african studies'], ['ethnic and racial studies '], ['[[nationalities papers'], ['turcica ', 'éditions klincksieck '], ['journal of the american oriental society '], ['the american journal of international law '], ['journal of world history '], ['journal of genocide research '], ['the british journal for the history of science ', '[[cambridge university press'], ['atlantic journal of communication '], ['middle eastern studies '], ['[[international studies quarterly'], ['international journal of middle east studies '], ['the journal of modern history '], ['journal for the history of astronomy ', 'science history publications ltd. '], ['cahiers du monde russe '], ['neurocirugía '], ['middle eastern studies '], ['urban development issues ']]",22278,Require autoconfirmed or confirmed access (no expiry set),229360,24 September 2001,BenBaker ,16644,30,2001-09-24,2001-09,2001
246,246,Vietnam,https://en.wikipedia.org/wiki/Vietnam,485,42,"['10.1355/sj16-1c', '10.17746/1563-0110.2018.46.3.003-021', '10.2112/jcoastres-d-16-00087.1', '10.2307/834104', '10.1016/j.scitotenv.2014.12.091', '10.1155/2014/528965', '10.1016/0022-5428(93)90038-q', '10.1127/zma/83/2001/59', '10.1016/s0304-4076(02)00161-6', '10.2307/2644255', '10.1355/sj11-1d', '10.1355/ae32-1c', '10.13140/2.1.5100.6249', '10.1038/s41467-020-19493-3', '10.1537/ase.070416', '10.1111/j.1365-3156.2005.01387.x', '10.3402/tellusa.v25i5.9694', '10.7152/bippa.v15i0.11537', '10.1080/10758216.2015.1083377', '10.1016/j.scitotenv.2006.09.010', '10.1111/j.1745-5871.2007.00487.x', '10.2307/3024603', '10.1016/j.proeng.2016.02.037', '10.2307/2761129', '10.1136/bmj.a137', '10.31235/osf.io/93fpa', '10.2307/2137774', '10.1525/as.2005.45.4.645', '10.2305/iucn.uk.2016-3.rlts.t45354985a95145107.en', '10.1016/j.proeng.2016.02.035', '10.1016/j.heliyon.2016.e00165', '10.1127/zma/77/1987/11', '10.2307/2645338', '10.1080/10871209.2018.1449038', '10.1596/1813-9450-2896', '10.1017/s0026749x00003590', '10.1038/scientificamerican0484-138', '10.1596/978-0-8213-7782-6', '10.1080/02549948.1976.11731121', '10.2307/3023970', '10.1355/cs22-2g', '19195125', None, None, None, '25585157', '24639878', None, '11372468', None, None, None, None, None, '33293507', None, '15807800', None, None, None, '17081593', None, None, None, None, '18566045', None, None, None, None, None, '27882357', '3564631', None, None, None, None, None, None, None, None, None, None, None, None, None, None, '3930020', None, None, None, None, None, None, None, '7723057', None, None, None, None, None, None, None, None, None, None, '2440905', None, None, None, None, None, '5114594', None, None, None, None, None, None, None, None, None, None]","[[' journal of social issues in southeast asia'], ['archaeology'], [' [[journal of coastal research'], ['  asian music'], [' [[science of the total environment'], [' journal of environmental and public health'], [' the columbia journal of world business'], [' zeitschrift für morphologie und anthropologie'], [' [[journal of econometrics'], ['  asian survey'], ['  sojourn'], [' southeast asian economies'], [' [[world bank'], ['nature communications'], [' anthropological science'], [' tropical medicine '], ['  tellus'], [' bulletin of the indo-pacific prehistory association'], [' [[problems of post-communism'], [' [[science of the total environment'], [' geographical research'], ['  far eastern survey'], [' procedia engineering'], ['  pacific affairs'], [' [[bmj'], ['pci archaeology '], [' population and development review'], ['[[asian survey', 'university of california press'], [' [[the iucn red list of threatened species'], [' procedia engineering'], [' heliyon'], [' zeitschrift für morphologie und anthropologie'], [' [[asian survey'], [' human dimensions of wildlife'], [' policy research working paper series'], [' [[modern asian studies'], [' scientific american'], [' [[world bank'], ['  monumenta serica'], ['  far eastern survey'], [' contemporary southeast asia']]",60,34,0,97,0,2,250,0.12371134020618557,0.07010309278350516,0.2,0.0865979381443299,0.0,0.2804123711340206,41,"['www.state.gov', 'www.moj.gov', 'xttm.agroviet.gov', 'teara.gov', 'www.mofa.gov', 'vietnamtourism.gov', 'www.mofa.gov', 'www.mofa.gov', 'agro.gov', '2009-2017.state.gov', 'www.usaid.gov', 'www.state.gov', 'minerals.usgs.gov', 'vbqppl.moj.gov', 'www.mofa.gov', '2009-2017.state.gov', 'luutru.gov', 'www.nea.gov', 'vbqppl.moj.gov', 'www.gso.gov', 'www.gov', 'files.eric.ed.gov', 'www.moj.gov', 'moj.gov', 'www.gov', 'dod.defense.gov', 'www.gso.gov', 'www.gov', 'vietnamtourism.gov', 'www.mofahcm.gov', 'www.gov', 'www.gso.gov', 'www.gso.gov', 'www.gso.gov', 'www.reuters.com', 'books.google.com', 'books.google.com', 'traveltips.usatoday.com', 'www.pwc.com', 'www.metalbulletin.com', 'www.oxfordscholarship.com', 'www.nytimes.com', 'www.thanhniennews.com', 'books.google.com', 'www.nytimes.com', 'www.vietnamonline.com', 'www.reuters.com', 'www.xinhuanet.com', 'www.nytimes.com', 'referenceworks.brillonline.com', 'www.scmp.com', 'www.vcsc.com', 'medium.com', 'books.google.com', 'worldview.stratfor.com', 'www.smentertainment.com', 'edition.cnn.com', 'www.thejakartapost.com', 'www.nytimes.com', 'www.popsci.com', 'thediplomat.com', 'gulfnews.com', 'books.google.com', 'news.google.com', 'books.google.com', 'www.techinasia.com', 'www.thanhniennews.com', 'www.agentorangerecord.com', 'www.duanemorris.com', 'books.google.com', 'english.chinamil.com', 'abc7news.com', 'www.formula1.com', 'www.ozy.com', 'books.google.com', 'news.com', 'socialistregister.com', 'www.vir.com', 'www.scmp.com', 'www.nytimes.com', 'www.evn.com', 'books.google.com', 'theaseanpost.com', 'www.indexmundi.com', 'www.history.com', 'books.google.com', 'www.universityworldnews.com', 'www.thecrimson.com', 'www.ecald.com', 'thediplomat.com', 'www.usatoday.com', 'theculturetrip.com', 'www.fourfourtwo.com', 'www.forbes.com', 'voices.yahoo.com', '2fwww.google.com', 'www.history.com', 'thediplomat.com', 'books.google.com', 'www.upi.com', 'asia.nikkei.com', 'www.nytimes.com', 'www.sbs.com', 'www.washingtonpost.com', 'www.bloomberg.com', 'economictimes.indiatimes.com', 'asia.nikkei.com', 'edition.cnn.com', 'oxfordbusinessgroup.com', 'thediplomat.com', 'www.indexmundi.com', 'books.google.com', 'www.historynet.com', 'www.saveur.com', 'thediplomat.com', 'asiatimes.com', 'www.economist.com', 'www.nytimes.com', 'scmp.com', 'matadornetwork.com', 'books.google.com', 'www.travelandleisure.com', 'allafrica.com', 'www.bbc.com', 'money.cnn.com', 'books.google.com', 'www.bbc.com', 'english.sina.com', 'www.nytimes.com', 'www.vir.com', 'www.bbc.com', 'treaties.un.org', 'en.nhandan.org', 'english.tapchicongsan.org', 'www.cuts-geneva.org', 'siteresources.worldbank.org', 'www.pri.org', 'thehuuvandan.org', 'data.worldbank.org', 'unesdoc.unesco.org', 'jahr.org', 'archives.the-monitor.org', 'www.popline.org', 'bbgv.org', 'www.imf.org', 'nationalinterest.org', 'mrlg.org', 'www.un.org', 'whc.unesco.org', 'www.tapchicongsan.org', 'data.worldbank.org', 'vietnamembassy-usa.org', 'whc.unesco.org', 'ich.unesco.org', 'population.un.org', 'fas.org', 'www.mhro.org', 'climatecentral.org', 'www.odi.org', 'data.worldbank.org', 'www.vn.undp.org', 'www.olympic.org', 'journals.openedition.org', 'data.worldbank.org', 'www.seaisi.org', 'www.unicef.org', 'www.odi.org', 'www.ohchr.org', 'www.seaaroundus.org', 'data.worldbank.org', 'vnsc.org', 'www.unesco.org', 'un-act.org', 'kyoto-seas.org', 'cpv.org', 'www.hoilhpn.org', 'hdr.undp.org', 'www.seafdec.org', 'data.worldbank.org', 'sggpnews.org', 'vietraleigh.org', 'www.unesco.org', 'www.riseprogramme.org', 'www.fwa.org', 'vietnam.unfpa.org', 'en.rsf.org', 'voxeu.org', 'data.worldbank.org', 'hdr.undp.org', 'washdata.org', 'data.worldbank.org', [' journal of social issues in southeast asia'], ['archaeology'], [' [[journal of coastal research'], ['  asian music'], [' [[science of the total environment'], [' journal of environmental and public health'], [' the columbia journal of world business'], [' zeitschrift für morphologie und anthropologie'], [' [[journal of econometrics'], ['  asian survey'], ['  sojourn'], [' southeast asian economies'], [' [[world bank'], ['nature communications'], [' anthropological science'], [' tropical medicine '], ['  tellus'], [' bulletin of the indo-pacific prehistory association'], [' [[problems of post-communism'], [' [[science of the total environment'], [' geographical research'], ['  far eastern survey'], [' procedia engineering'], ['  pacific affairs'], [' [[bmj'], ['pci archaeology '], [' population and development review'], ['[[asian survey', 'university of california press'], [' [[the iucn red list of threatened species'], [' procedia engineering'], [' heliyon'], [' zeitschrift für morphologie und anthropologie'], [' [[asian survey'], [' human dimensions of wildlife'], [' policy research working paper series'], [' [[modern asian studies'], [' scientific american'], [' [[world bank'], ['  monumenta serica'], ['  far eastern survey'], [' contemporary southeast asia']]",202354,Require administrator access (no expiry set),310552,27 March 2001,TimShell ,10581,11,2001-03-27,2001-03,2001
247,247,Griko people,https://en.wikipedia.org/wiki/Griko_people,92,0,[],[],0,1,0,16,0,0,76,0.0,0.010869565217391304,0.17391304347826086,0.0,0.0,0.010869565217391304,0,"['www.greciasalentina.gov', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.com', 'books.google.com', 'books.google.com', 'www.amazon.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'greece.greekreporter.com', 'books.google.com', 'books.google.com', 'books.google.com']",30804808,Allow all users (no expiry set),81658,9 February 2011,Runselit ,365,3,2011-02-09,2011-02,2011
248,248,Mangalore,https://en.wikipedia.org/wiki/Mangalore,410,1,"[None, None, 'pdfw.mr']",[['mangalore refinery and petrochemicals ']],5,18,0,299,0,0,87,0.012195121951219513,0.04390243902439024,0.7292682926829268,0.0024390243902439024,0.0,0.05853658536585366,1,"['censuskarnataka.gov', 'www.mangalorecity.gov', 'imdpune.gov', 'imdpune.gov', 'censusindia.gov', 'imdpune.gov', 'www.mangalorecity.gov', 'www.censusindia.gov', 'censusindia.gov', 'customsmangalore.gov', 'www.mangalorecity.gov', 'gcmd.nasa.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'imdpune.gov', 'www.mangalorecity.gov', 'www.imdbangalore.gov', 'cgwb.gov', 'www.thehindu.com', 'www.daijiworld.com', 'www.thehindu.com', 'www.daijiworld.com', 'www.thehindu.com', 'www.mapsofindia.com', 'www.thehindu.com', 'www.thehindu.com', 'articles.timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.w3newspapers.com', 'www.business-standard.com', 'www.deccanherald.com', 'timesofindia.indiatimes.com', 'www.hindu.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', '2fmangalorean.com', 'www.thehindu.com', 'books.google.com', 'www.thehindubusinessline.com', 'www.deccanherald.com', 'www.thehindubusinessline.com', 'www.thehindu.com', 'www.deccanherald.com', 'www.thehindu.com', 'www.thehindu.com', 'www.daijiworld.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.indiacom.com', 'v4news.com', 'www.dnaindia.com', 'articles.timesofindia.indiatimes.com', 'www.thehindu.com', 'www.daijiworld.com', 'www.konkanrailway.com', 'www.hindu.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.deccanherald.com', 'www.thehindu.com', 'www.thehindu.com', 'mangalorean.com', 'www.thehindu.com', 'www.bellevision.com', 'www.deccanherald.com', 'www.thehindu.com', 'weather-and-climate.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.deccanherald.com', 'www.hindu.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.com', 'www.thehindu.com', 'www.thehindu.com', 'cincinnatitemple.com', 'www.daijiworld.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.deccanherald.com', 'www.mangalorean.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.daijiworld.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'profit.ndtv.com', 'timesofindia.indiatimes.com', 'content-www.cricinfo.com', 'www.pilikula.com', 'www.thehindubusinessline.com', 'english.mathrubhumi.com', 'www.scdccbank.com', 'www.thehindubusinessline.com', 'www.thehindu.com', 'hindu.com', 'www.konkanworld.com', 'www.weatherbase.com', 'www.thehindu.com', 'www.mangaloretoday.com', 'www.thehindubusinessline.com', 'www.thehindu.com', 'www.thehindu.com', 'www.deccanherald.com', 'www.business-standard.com', 'timesofindia.indiatimes.com', 'bangaloremirror.indiatimes.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'www.deccanherald.com', 'www.deccanchronicle.com', 'www.hindu.com', 'www.thehindu.com', 'www.hindu.com', 'www.corpbank.com', 'www.deccanherald.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'economictimes.indiatimes.com', 'archive.deccanherald.com', 'www.thehindu.com', 'www.deccanherald.com', 'books.google.com', 'archive.deccanherald.com', 'archive.deccanherald.com', 'www.thehindu.com', 'content-www.cricinfo.com', '2fwww.daijiworld.com', 'www.thehindu.com', 'www.deccanherald.com', 'www.daijiworld.com', 'www.daijiworld.com', 'books.google.com', 'www.deccanherald.com', 'vijayabank.com', 'timesofindia.indiatimes.com', 'www.hindu.com', 'www.thehindu.com', 'www.daijiworld.com', 'www.heraldmalaysia.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.thehindubusinessline.com', 'www.karnatakabank.com', 'www.deccanchronicle.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.daijiworld.com', 'www.thehindu.com', 'www.epapermathrubhumi.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'www.deccanherald.com', 'www.thehindu.com', 'coastaldigest.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.thehindu.com', 'karnataka.com', 'www.hindu.com', 'books.google.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.daijiworld.com', 'www.daijiworld.com', 'www.thehindu.com', 'www.thehindu.com', 'www.business-standard.com', 'mangalorean.com', 'www.deccanherald.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.daijiworld.com', 'www.thehindubusinessline.com', 'www.hindu.com', 'www.hindu.com', 'www.thehindu.com', 'www.business-standard.com', 'www.daijiworld.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehindu.com', 'www.daijiworld.com', 'www.thehindu.com', 'www.daijiworld.com', 'economictimes.indiatimes.com', 'www.daijiworld.com', 'www.deccanherald.com', 'www.business-standard.com', 'www.thehindubusinessline.com', 'timesofindia.indiatimes.com', 'www.deccanherald.com', 'www.deccanherald.com', 'www.outlookindia.com', 'www.thehindubusinessline.com', 'www.thehindu.com', 'www.business-standard.com', 'www.sportskeeda.com', 'www.thehindu.com', 'books.google.com', 'www.daijiworld.com', 'www.karnatakachess.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'www.geographicus.com', 'articles.timesofindia.indiatimes.com', 'www.daijiworld.com', 'www.daijiworld.com', 'www.deccanherald.com', 'www.thehindu.com', 'www.deccanherald.com', 'www.thehindu.com', 'www.karnataka.com', 'indianexpress.com', 'www.timesnownews.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.thehindu.com', 'www.financialexpress.com', 'www.deccanherald.com', 'timesofindia.indiatimes.com', 'www.daijiworld.com', 'www.medianewsline.com', 'timesofindia.indiatimes.com', 'www.thehindubusinessline.com', 'www.deccanherald.com', '2fwww.daijiworld.com', 'timesofindia.indiatimes.com', 'www.deccanherald.com', 'books.google.com', 'www.thenewsminute.com', 'm.timesofindia.com', 'www.hindu.com', 'canaratv.com', 'www.deccanherald.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.thehindu.com', 'www.daijiworld.com', 'www.nammakudlanews.com', 'www.thenewsminute.com', 'timesofindia.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.thehindu.com', 'www.thehindu.com', 'www.daijiworld.com', 'www.fallingrain.com', 'timesofindia.indiatimes.com', 'www.educationobserver.com', 'www.daijiworld.com', 'www.hindu.com', 'books.google.com', 'archive.deccanherald.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.thehindubusinessline.com', 'content-www.cricinfo.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehindu.com', '2fwww.karavaliutsav.com', 'www.thehindu.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'www.thehindu.com', 'www.epapermathrubhumi.com', 'www.hindu.com', 'www.hindu.com', 'www.thehindubusinessline.com', 'economictimes.indiatimes.com', 'books.google.com', 'www.konkanworld.com', 'www.hindu.com', 'www.thehindu.com', 'www.business-standard.com', 'timesofindia.indiatimes.com', 'content-usa.cricinfo.com', 'www.daijiworld.com', 'www.thehindu.com', 'www.hindu.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehindu.com', 'www.epapersland.com', 'www.deccanherald.com', 'www.mangalorechemicals.com', 'timesofindia.com', 'books.google.com', 'www.kptcl.com', 'www.deccanherald.com', 'economictimes.indiatimes.com', 'www.hindu.com', 'indianexpress.com', 'whc.unesco.org', 'www.commonlii.org', 'www.nio.org', 'www.nhai.org', '2fwww.tertullian.org', ['mangalore refinery and petrochemicals ']]",308293,Require administrator access (no expiry set),188436,31 August 2003,Pradeep bt ,8982,3,2003-08-31,2003-08,2003
249,249,Mali,https://en.wikipedia.org/wiki/Mali,175,3,"['10.2307/634762', '10.1093/biosci/bix014', '10.1038/s41467-020-19493-3', None, '28608869', '33293507', None, '5451287', '7723057']","[['the geographical journal'], ['bioscience'], ['nature communications']]",36,10,0,51,0,5,70,0.2057142857142857,0.05714285714285714,0.2914285714285714,0.017142857142857144,0.0,0.28,3,"['www.cia.gov', 'www.usaid.gov', 'www.cia.gov', 'lcweb2.loc.gov', 'www.matcl.gov', '2009-2017.state.gov', 'instat.gov', 'www.cia.gov', 'www.usaid.gov', 'state.gov', 'fr.allafrica.com', 'foreignpolicy.com', 'www.indexmundi.com', 'www.kirasalak.com', 'books.google.com', 'www.sedar.com', 'www.britannica.com', 'news.nationalgeographic.com', 'www.bbc.com', 'www.aa.com', 'malijet.com', 'www.aljazeera.com', 'www.aljazeera.com', 'edition.cnn.com', 'dhsprogram.com', 'www.nytimes.com', 'www.france24.com', 'www.best-country.com', 'report.com', 'abcnews.go.com', 'www.bbc.com', '.com', 'www.reuters.com', 'www.aljazeera.com', 'www.theglobeandmail.com', 'www.google.com', 'www.aljazeera.com', 'www.sfgate.com', 'www.nytimes.com', 'threadster.com', 'www.usatoday.com', 'www.nytimes.com', 'www.fivb.com', 'blog.namsor.com', 'africanews.com', 'www.aljazeera.com', 'books.google.com', 'www.africanews.com', 'www.aljazeera.com', 'www.news24.com', 'books.google.com', 'www.theglobeandmail.com', 'www.ohada.com', 'www.indexmundi.com', 'books.google.com', 'www.bbc.com', 'www.ibtimes.com', 'books.google.com', 'books.google.com', 'africabasket.com', 'aglobalworld.com', 'world-nuclear.org', 'africanarguments.org', 'www.imf.org', 'www.hdcentre.org', 'www.hdcentre.org', 'blackpast.org', 'wise-uranium.org', 'hdr.undp.org', 'www.undp.org', 'data.un.org', 'www.ictj.org', 'en.puic.org', 'www.instat-mali.org', 'news.un.org', 'www.thenewhumanitarian.org', 'www.nonviolent-conflict.org', 'www.wto.org', 'promundoglobal.org', 'www.pewforum.org', 'minusma.unmissions.org', 'www.instat-mali.org', 'ambamali-jp.org', 'www.nonviolent-conflict.org', 'minusma.unmissions.org', 'www.nationalgeographic.org', 'data.worldbank.org', 'www.nonviolent-conflict.org', 'www.worldbank.org', 'www.omct.org', 'hdr.undp.org', 'unpan1.un.org', 'datatopics.worldbank.org', 'www.hrw.org', 'hdr.undp.org', 'www.hrw.org', 'www.impatientoptimists.org', ['the geographical journal'], ['bioscience'], ['nature communications']]",19127,Require administrator access (no expiry set),130384,28 September 2001,Koyaanis Qatsi ,5112,30,2001-09-28,2001-09,2001
250,250,Culture of Europe,https://en.wikipedia.org/wiki/Culture_of_Europe,36,0,[],[],3,0,0,3,0,0,30,0.08333333333333333,0.0,0.08333333333333333,0.0,0.0,0.08333333333333333,0,"['www.journeywonders.com', 'sciendo.com', 'europeword.com', 'www.pewforum.org', 'pewforum.org', 'pewforum.org']",1256013,Allow all users (no expiry set),63072,8 December 2004,Thewayforward ,2300,2,2004-12-08,2004-12,2004
251,251,Ibiza,https://en.wikipedia.org/wiki/Ibiza,55,1,"['10.1353/pgn.2013.0016', None, None]",[['parergon']],6,0,0,19,0,3,26,0.10909090909090909,0.0,0.34545454545454546,0.01818181818181818,0.0,0.12727272727272726,1,"['www.billboard.com', 'www.petitfute.com', 'www.healingibiza.com', 'www.liveibiza.com', 'www.vipealo.com', 'ibizaphoto.blogspot.com', 'www.bbc.com', 'www.vice.com', 'www.ibizatraveller.com', 'ibizaphoto.blogspot.com', 'www.directferries.com', 'gointothestory.blcklst.com', 'irenedeandres.com', 'www.resortsinspain.com', 'ibizaphoto.blogspot.com', 'books.google.com', 'liveibiza.com', 'bbs.clubplanet.com', 'www.weather-atlas.com', 'whc.unesco.org', 'tvtropes.org', 'seatemperature.org', 'www.seatemperature.org', 'www.travelntourism.org', 'whc.unesco.org', ['parergon']]",63624,Allow all users (no expiry set),46245,23 July 2002,Perique des Palottes ,3072,1,2002-07-23,2002-07,2002
252,252,Madrid,https://en.wikipedia.org/wiki/Madrid,232,8,"['10.14198/ingeo2016.66.03', '10.14483/22487638.6249', '10.4000/argonauta.4257', '10.1017/s0963926800000808', '10.4067/s0718-93032016000200013', '10.1080/14649360701633212', '10.1080/01441640802383214', '10.1002/kpm.346', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None]","[['investigaciones geográficas'], ['tecnura', '[[francisco josé de caldas district university'], ['el argonauta español'], ['[[urban history'], ['boletín de filología'], ['[[taylor ', 'social '], ['transport reviews'], ['knowledge and process management ']]",11,0,0,82,0,2,129,0.04741379310344827,0.0,0.35344827586206895,0.034482758620689655,0.0,0.08189655172413793,8,"['elpais.com', 'www.alimente.elconfidencial.com', 'www.audiovisual451.com', 'global.britannica.com', 'www.nytimes.com', 'books.google.com', 'www.lavanguardia.com', 'timeout.com', 'books.google.com', 'www.lavanguardia.com', 'www.demographia.com', 'variety.com', 'forbes.com', 'historialia.com', 'mercedesbenzfashionweekmadrid.com', 'www.reuters.com', 'www.libremercado.com', 'www.lavanguardia.com', 'www.esmadrid.com', 'www.nytimes.com', 'nileguide.com', 'elpais.com', 'escenacontemporanea.com', 'sincro.com', 'gomadrid.com', 'www.lasexta.com', 'elpais.com', 'elpais.com', 'www.madridorgullo.com', 'www.citymayors.com', 'elpais.com', 'elmadridmedieval.jmcastellanos.com', 'www.broadbandtvnews.com', 'www.airport-technology.com', 'www.elespanol.com', 'elpais.com', 'elpais.com', 'elpais.com', 'www.economiademadrid.com', 'www.madrid-destino.com', 'elpais.com', 'www.nytimes.com', 'www.highbeam.com', 'www.easyexpat.com', 'www.mastercard.com', 'elpais.com', 'www.lavanguardia.com', 'www.easyexpat.com', 'www.alimente.elconfidencial.com', 'www.demographia.com', 'www.ukmediacentre.pwc.com', 'books.google.com', 'indigoguide.com', 'noticias.juridicas.com', 'www.timeout.com', 'whatmadrid.com', 'elpais.com', 'books.google.com', 'notesfrommadrid.com', 'inhabitat.com', 'books.google.com', 'www.goal.com', 'elpais.com', 'www.madrid-traveller.com', 'elpais.com', 'en.momondo.com', 'www.redforesta.com', 'www.thejakartapost.com', 'www.audiovisual451.com', 'elpais.com', 'www.highbeam.com', 'elpais.com', 'www.bbc.com', 'elpais.com', 'www.timeout.com', 'www.citylab.com', 'cronicaglobal.elespanol.com', 'elpais.com', 'cincodias.elpais.com', 'www.madridorgullo.com', 'www.lavanguardia.com', 'cnn.com', 'hdi.globaldatalab.org', 'www.un.org', 'www.madrid.org', 'books.openedition.org', 'www.madrid.org', 'www.oschamartin.org', 'www.museothyssen.org', 'www.madrid.org', 'secforestales.org', 'www.madrid.org', 'www.tiemposmodernos.org', ['investigaciones geográficas'], ['tecnura', '[[francisco josé de caldas district university'], ['el argonauta español'], ['[[urban history'], ['boletín de filología'], ['[[taylor ', 'social '], ['transport reviews'], ['knowledge and process management ']]",41188263,Require administrator access (no expiry set),210126,18 December 2001,147.83.41.xxx ,10626,12,2001-12-18,2001-12,2001
253,253,Greek Cypriots,https://en.wikipedia.org/wiki/Greek_Cypriots,19,4,"['10.21773/boun.25.2.6', '10.1038/nature23310', '10.1038/s41598-017-01802-4', '10.1371/journal.pone.0179474', None, '28783727', '28512355', '28622394', None, '5565772', '5434004', '5473566']","[['bogazici journal '], ['[[nature '], ['[[scientific reports'], ['[[plos one']]",1,5,0,4,0,0,5,0.05263157894736842,0.2631578947368421,0.21052631578947367,0.21052631578947367,0.0,0.5263157894736842,4,"['lcweb2.loc.gov', 'www.cyprus.gov', 'www.cyprus.gov', 'www.cystat.gov', 'www.cyprus.gov', 'ςww.apotipomata.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.cnewa.org', ['bogazici journal '], ['[[nature '], ['[[scientific reports'], ['[[plos one']]",1210883,Allow all users (no expiry set),28373,26 November 2004,66.25.176.71 ,838,15,2004-11-26,2004-11,2004
254,254,Kosovo,https://en.wikipedia.org/wiki/Kosovo,275,6,"['10.1163/187633009x411485', '10.1093/biosci/bix014', '10.5771/0506-7286-1999-3-422', '10.1080/13602000903411366', '10.1023/a:1025397128633', '10.1038/s41467-020-19493-3', None, '28608869', None, None, None, '33293507', None, '5451287', None, None, None, '7723057']","[['east central europe'], ['bioscience'], ['verfassung in recht und übersee'], ['journal of muslim minority affairs'], ['international journal of politics'], ['nature communications']]",59,12,0,77,0,3,118,0.21454545454545454,0.04363636363636364,0.28,0.02181818181818182,0.0,0.28,6,"['www.instat.gov', 'pdf.usaid.gov', 'www.serbia.sr.gov', 'pdf.usaid.gov', 'www.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'buyusa.gov', 'www.sam.gov', 'parlament.gov', 'www.srbija.gov', 'www.dw.com', 'freethoughtreport.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'uk.reuters.com', 'www.jpost.com', 'travel.nytimes.com', 'webcache.googleusercontent.com', 'www.foreignaffairs.com', 'books.google.com', 'books.google.com', 'rebibneenun.blogdetik.com', 'www.fiba.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'balkaninsight.com', 'www.itg-rks.com', 'books.google.com', 'books.google.com', 'www.eonline.com', 'books.google.com', 'www.hollywoodreporter.com', 'books.google.com', 'rio2016.com', 'prishtinainsight.com', 'books.google.com', 'rs.n1info.com', 'www.alb-net.com', 'www.hollywoodreporter.com', 'www.podravka.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'adnkronos.com', 'prishtinainsight.com', 'setimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'setimes.com', 'rs.n1info.com', 'books.google.com', 'books.google.com', 'kosovareport.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'webcache.googleusercontent.com', 'books.google.com', 'www.economist.com', 'www.dokufest.com', 'content.time.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'www.trainkos.com', 'www.france24.com', 'books.google.com', 'worldpopulationreview.com', 'books.google.com', 'www.ft.com', 'kosovapress.com', 'www.britannica.com', 'www.setimes.com', 'books.google.com', 'heritage.sense-agency.com', 'kosovotwopointzero.com', 'balkaninsight.com', 'www.voanews.com', 'www.eciks.org', 'icty.org', 'esiweb.org', 'www.hrw.org', 'mksf-ks.org', 'www.mti-ks.org', 'www.unesco.org', 'constituteproject.org', 'mmph-rks.org', 'unstats.un.org', 'constituteproject.org', 'olympic.org', 'www.unhcr.org', 'whc.unesco.org', 'www.kosovomemorybook.org', 'visionofhumanity.org', 'kcr-ks.org', 'www.unhcr.org', 'icty.org', 'icty.org', 'www.eciks.org', 'www.hrw.org', 'icty.org', 'www.kosovo-mining.org', 'internal-displacement.org', 'constituteproject.org', 'web.worldbank.org', 'www.cpa.org', 'www.imf.org', 'www.osce.org', 'www.mkrs-ks.org', 'www.imf.org', 'euinkosovo.org', 'qkuk.org', 'data.worldbank.org', 'euinkosovo.org', 'publicinternationallaw.org', 'www.kosovo-mining.org', 'www.kosovo-eicc.org', 'www.esiweb.org', 'internal-displacement.org', 'www.irex.org', 'imf.org', 'icj-cij.org', 'whc.unesco.org', 'www.osce.org', 'whc.unesco.org', 'www.icj-cij.org', 'www.hrw.org', 'mksf-ks.org', 'siteresources.worldbank.org', 'dissidentvoice.org', 'www.osce.org', 'www.prishtina-komuna.org', 'www.osce.org', 'www.osce.org', 'hdr.undp.org', 'msh-ks.org', 'constituteproject.org', ['east central europe'], ['bioscience'], ['verfassung in recht und übersee'], ['journal of muslim minority affairs'], ['international journal of politics'], ['nature communications']]",17391,Require administrator access (no expiry set),225096,15 December 2001,Hagedis ,13445,23,2001-12-15,2001-12,2001
255,255,"Tarsus, Mersin","https://en.wikipedia.org/wiki/Tarsus,_Mersin",23,3,"['10.1163/1877837292x00105', '10.2307/596170', None, None, None, None]","[[' oriens '], [' journal of the american oriental society ']]",1,0,0,2,0,0,17,0.043478260869565216,0.0,0.08695652173913043,0.13043478260869565,0.0,0.17391304347826086,2,"['books.google.com', 'www.jewishencyclopedia.com', 'www.wdl.org', [' oriens '], [' journal of the american oriental society ']]",871713,Allow all users (no expiry set),36098,1 August 2004,Yak ,748,0,2004-08-01,2004-08,2004
256,256,Altai people,https://en.wikipedia.org/wiki/Altai_people,40,11,"['10.1038/s41586-018-0094-2', '10.1163/22105832-00702005', '10.1017/ehs.2020.11', '10.1017/ehs.2020.4', None, '10.1016/j.ara.2020.100177', '10.1080/1361736042000245295', '10.1016/j.ajhg.2011.12.014', '10.4000/emscat.2444', '10.1163/22105018-12340089', '10.2753/aae1061-1959450303', '10.1038/srep20768', '29743675', None, None, None, None, None, None, '22281367', None, None, None, '26865217', None, None, None, None, None, None, None, '3276666', None, None, None, '4750364']","[['[[nature ', '[[nature research'], ['language dynamics and change ', '[[brill publishers'], ['evolutionary human sciences ', '[[cambridge university press'], ['evolutionary human sciences ', '[[cambridge university press'], ['журнал социологии и социальной антропологии [journal of sociology and social anthropology'], ['archaeological research in asia ', '[[elsevier'], ['sibirica '], ['the american journal of human genetics'], ['études mongoles et sibériennes'], ['inner asia ', '[[brill publishers'], ['anthropology '], ['scientific reports']]",0,0,0,12,0,0,16,0.0,0.0,0.3,0.275,0.0,0.275,12,"['books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.pressreader.com', 'books.google.com', 'global.oup.com', 'books.google.com', 'www.endangeredlanguages.com', 'books.google.com', ['[[nature ', '[[nature research'], ['language dynamics and change ', '[[brill publishers'], ['evolutionary human sciences ', '[[cambridge university press'], ['evolutionary human sciences ', '[[cambridge university press'], ['журнал социологии и социальной антропологии [journal of sociology and social anthropology'], ['archaeological research in asia ', '[[elsevier'], ['sibirica '], ['the american journal of human genetics'], ['études mongoles et sibériennes'], ['inner asia ', '[[brill publishers'], ['anthropology '], ['scientific reports']]",4878363,Allow all users (no expiry set),33435,24 April 2006,Imz ,421,6,2006-04-24,2006-04,2006
257,257,Dogras,https://en.wikipedia.org/wiki/Dogras,13,0,[],[],1,2,0,7,0,0,3,0.07692307692307693,0.15384615384615385,0.5384615384615384,0.0,0.0,0.23076923076923078,0,"['censusindia.gov', 'jammutourism.gov', 'duggartimes.com', 'www.tribuneindia.com', 'books.google.com', 'webindia123.com', 'books.google.com', 'www.tribuneindia.com', 'books.google.com', 'globalsecurity.org']",1823707,Allow all users (no expiry set),17958,1 May 2005,Rl ,1576,9,2005-05-01,2005-05,2005
258,258,Prague,https://en.wikipedia.org/wiki/Prague,149,1,[],[],12,2,0,49,0,0,85,0.08053691275167785,0.013422818791946308,0.3288590604026846,0.006711409395973154,0.0,0.10067114093959731,0,"['ftp.atdd.noaa.gov', 'www.miamidade.gov', 'abcprague.com', 'mobilityexchange.mercer.com', 'www.praguepost.com', 'books.google.com', 'tripadvisor.com', 'books.google.com', 'books.google.com', 'www.chicagosistercities.com', 'czech-transport.com', 'books.google.com', 'books.google.com', 'praguemonitor.com', 'mobilityexchange.mercer.com', 'www.pragueexperience.com', 'www.travelmath.com', 'demographia.com', 'worldatlas.com', 'worldatlas.com', 'praguestudios.com', 'www.infoplease.com', 'www.theartnewspaper.com', 'www.myczechrepublic.com', 'www.architecturaldigest.com', 'piscaindex.com', 'portal.com', 'books.google.com', 'eiuresources.com', 'www.worldinfozone.com', 'nakedtourguideprague.com', 'www.praguepost.com', 'www.gamesbids.com', 'www.architecturaldigest.com', 'www.innovation-cities.com', 'www.praguepost.com', 'books.google.com', 'railwaytechnology.com', 'www.newprague.com', 'www.praguepost.com', 'books.google.com', 'www.worldinfozone.com', 'praguesummer.com', 'www.weatherbase.com', 'cs-magazin.com', 'euobserver.com', 'www.weather-atlas.com', 'gamesbids.com', 'thediplomat.com', 'books.google.com', 'www.infoplease.com', 'www.phoenixsistercities.org', 'www.iajgsjewishcemeteryproject.org', 'brrp.org', 'www.everything2.org', 'cityofpragueok.org', 'hdi.globaldatalab.org', 'tshaonline.org', 'libmma.contentdm.oclc.org', 'www.hebrewbooks.org', 'www.peoplesworld.org', 'wfdf.org', 'www.jewishvirtuallibrary.org']",23844,Require administrator access (no expiry set),148315,6 November 2001,WojPob ,6096,21,2001-11-06,2001-11,2001
259,259,Culture of Spain,https://en.wikipedia.org/wiki/Culture_of_Spain,17,2,"['10.1080/10286632.2018.1514036', '10.1057/9781137531070.0010', None, None, None, None]","[['international journal of cultural policy'], ['brill']]",2,0,0,2,0,0,11,0.11764705882352941,0.0,0.11764705882352941,0.11764705882352941,0.0,0.23529411764705882,2,"['ethnologue.com', 'www.dw.com', 'www.realinstitutoelcano.org', 'whc.unesco.org', ['international journal of cultural policy'], ['brill']]",1010051,Allow all users (no expiry set),33291,23 September 2004,Taxman ,2162,1,2004-09-23,2004-09,2004
260,260,Jharkhand,https://en.wikipedia.org/wiki/Jharkhand,138,2,"['10.11588/xarep.00000510', '10.1007/s00223-005-0233-2', None, '15895280', None, None]","[['man in environment'], ['calcified tissue international']]",13,11,0,71,0,0,41,0.09420289855072464,0.07971014492753623,0.5144927536231884,0.014492753623188406,0.0,0.18840579710144928,2,"['census.gov', 'www.censusindia.gov', 'censusindia.gov', 'jharkhandtourism.gov', 'www.jharkhand.gov', 'www.wii.gov', 'www.jharkhand.gov', 'www.censusindia.gov', 'censusindia.gov', 'www.jharkhand.gov', 'censusindia.gov', 'www.atimes.com', 'www.dailypioneer.com', 'www.dailypioneer.com', 'www.telegraphindia.com', 'educationforallinindia.com', 'www.telegraphindia.com', 'indianvagabond.com', 'www.telegraphindia.com', 'articles.timesofindia.indiatimes.com', 'mapsofindia.com', 'www.telegraphindia.com', 'india.com', 'tourism.webindia123.com', 'economictimes.indiatimes.com', 'www.dailypioneer.com', 'www.dailypioneer.com', 'www.laureus.com', 'www.disabled-world.com', 'business.mapsofindia.com', 'www.telegraphindia.com', 'books.google.com', 'www.globalpolitician.com', 'books.google.com', 'www.ndtv.com', 'www.thehindu.com', 'www.southasiaarchive.com', 'www.mapsofindia.com', 'www.telegraphindia.com', 'www.telegraphindia.com', 'jharkhandstatenews.com', 'www.telegraphindia.com', 'timesofindia.indiatimes.com', 'tatamemorialcentre.com', 'news.webindia123.com', 'www.thehindu.com', 'www.uniindia.com', 'traveljharkhand.com', 'business.rediff.com', 'books.google.com', 'www.telegraphindia.com', 'india.com', 'hindustantimes.com', 'ndtv.com', 'www.hindustantimes.com', 'nyoooz.com', 'www.moneycontrol.com', 'www.business-standard.com', 'www.outlookindia.com', 'prabhatkhabar.com', 'books.google.com', 'www.telegraphindia.com', 'roadtraffic-technology.com', 'www.telegraphindia.com', 'www.dailypioneer.com', 'mdaily.bhaskar.com', 'books.google.com', 'www.nytimes.com', 'www.thehindu.com', 'www.hindustantimes.com', 'books.google.com', 'www.dailypioneer.com', 'www.newindianexpress.com', 'books.google.com', 'www.telegraphindia.com', 'www.telegraphindia.com', 'm.jagranjosh.com', 'books.google.com', 'articles.timesofindia.indiatimes.com', 'www.telegraphindia.com', 'www.business-standard.com', 'timesofindia.indiatimes.com', 'gandhiserve.org', 'sa.indiaenvironmentportal.org', 'www.prsindia.org', 'www.ibef.org', 'www.nhai.org', 'www.gandhimedia.org', 'www.ibef.org', 'en.climate-data.org', 'www.mkgandhi-sarvodaya.org', 'www.nfhsindia.org', 'www.in.undp.org', 'www.aicc.org', 'www.asiranchi.org', ['man in environment'], ['calcified tissue international']]",197225,Allow all users (no expiry set),115540,16 March 2003,202.141.140.133 ,5554,30,2003-03-16,2003-03,2003
261,261,Bulgarians,https://en.wikipedia.org/wiki/Bulgarians,177,3,"['10.1556/aorient.58.2005.1.1', '0584-9888/2010/0584-98881047055k.pdf', '10.1371/journal.pone.0135820', None, None, '26332464', None, None, '4558026']","[['acta orientalia academiae scientiarum hungaricae '], ['зборник радова византолошког института'], ['plos one ']]",5,7,0,75,0,0,87,0.02824858757062147,0.03954802259887006,0.423728813559322,0.01694915254237288,0.0,0.0847457627118644,3,"['factfinder.census.gov', 'abs.gov', 'www.stat.gov', 'aba.gov', 'ons.gov', 'cystat.gov', 'ukrcensus.gov', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'macedonia.kroraina.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'fcbarcelona.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.kroraina.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.protobulgarians.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thepoultrysite.com', 'books.google.com', 'www.maritsa.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'kroraina.com', 'books.google.com', 'etnoxata.com', 'books.google.com', 'www.ceeol.com', 'books.google.com', 'books.google.com', 'kroraina.com', 'books.google.com', 'www.milliyet.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.ethnologue.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'kroraina.com', 'books.google.com', 'www.keepeek.com', 'tangrabg.files.wordpress.com', 'kroraina.com', 's7.hostingkartinok.com', 'promacedonia.org', 'promacedonia.org', 'pop-stat.mashke.org', 'bkks.org', 'promacedonia.org', ['acta orientalia academiae scientiarum hungaricae '], ['зборник радова византолошког института'], ['plos one ']]",151876,Allow all users (no expiry set),113991,26 November 2002,195.170.20.8 ,6269,10,2002-11-26,2002-11,2002
262,262,"Punjab, India","https://en.wikipedia.org/wiki/Punjab,_India",196,1,"['10.2752/147800409x466254', None, None]",[['cultural and social history']],11,21,0,103,0,1,60,0.05612244897959184,0.10714285714285714,0.5255102040816326,0.00510204081632653,0.0,0.1683673469387755,1,"['ftp.atdd.noaa.gov', 'mhrd.gov', 'www.indianrailways.gov', 'data.gov', 'imdpune.gov', 'censusindia.gov', 'www.mospi.gov', 'census.gov', 'censusindia.gov', 'agriexchange.apeda.gov', 'punjabgovt.gov', 'censusindia.gov', 'www.censusindia.gov', 'pbplanning.gov', 'imdpune.gov', 'punjab.gov', 'censusindia.gov', 'agriexchange.apeda.gov', 'www.nfsm.gov', 'censusindia.gov', 'censusindia.gov', 'zeenews.india.com', 'www.huffingtonpost.com', 'food.ndtv.com', 'www.dayandnightnews.com', 'indianexpress.com', 'books.google.com', 'www.tribuneindia.com', 'www.afaqs.com', 'www.kamloopsthisweek.com', 'www.tribuneindia.com', 'www.tribuneindia.com', 'www.discoveredindia.com', 'timesofindia.indiatimes.com', 'www.business-standard.com', 'www.bollywoodlife.com', 'zeenews.india.com', 'www.news18.com', 'timesofindia.indiatimes.com', 'www.hindustantimes.com', 'food.ndtv.com', 'www.thehindu.com', 'www.hindustantimes.com', 'www.radioandmusic.com', 'www.appeal-democrat.com', 'www.britannica.com', 'www.tribuneindia.com', 'www.nytimes.com', 'timesofindia.indiatimes.com', 'www.tribuneindia.com', 'timesofindia.indiatimes.com', 'www.telegraphindia.com', 'books.google.com', 'mapsofindia.com', 'economictimes.indiatimes.com', 'www.ibtimes.com', 'www.hindustantimes.com', 'www.thehindu.com', 'www.thehindubusinessline.com', 'www.hindustantimes.com', 'www.hindustantimes.com', 'www.livemint.com', 'www.philly.com', 'food.ndtv.com', 'www.newindianexpress.com', 'indianexpress.com', 'books.google.com', 'indianexpress.com', 'archive.indiaspend.com', 'www.tribuneindia.com', 'punjabilok.com', 'www.discoveredindia.com', 'www.discoveredindia.com', 'books.google.com', 'books.google.com', 'tns.thenews.com', 'www.globalpunjabtv.com', 'www.brantnews.com', 'www.firstpost.com', 'books.google.com', 'www.statista.com', 'books.google.com', 'books.google.com', 'www.hindustantimes.com', 'books.google.com', 'www.bbc.com', 'www.business-standard.com', 'www.indiatvnews.com', 'indianexpress.com', 'www.indiatvnews.com', 'www.dailytimes.com', 'timesofindia.indiatimes.com', 'archive.indianexpress.com', 'www.thefridaytimes.com', 'ptinews.com', 'zeenews.india.com', 'www.ebc-india.com', 'tribune.com', 'www.indiantelevision.com', 'timesofindia.indiatimes.com', 'nba.com', 'www.indiantelevision.com', 'www.tribuneindia.com', 'www.google.com', 'economictimes.indiatimes.com', 'www.wsj.com', 'economictimes.indiatimes.com', 'www.deccanherald.com', 'www.britannica.com', 'books.google.com', 'www.exoticindiaart.com', 'www.mapsofindia.com', 'www.newindianexpress.com', 'www.desiblitz.com', 'www.indiantelevision.com', 'books.google.com', 'www.britannica.com', 'www.asiantribune.com', 'www.hindustantimes.com', 'www.bhaskar.com', 'books.google.com', 'www.hindustantimes.com', 'www.thehindu.com', 'books.google.com', 'cpasindia.org', 'www.filmfed.org', 'www.filmfed.org', 'rbidocs.rbi.org', 'hdi.globaldatalab.org', 'www.circleofblue.org', 'bhangra.org', 'ich.unesco.org', 'www.gutenberg.org', 'www.gutenberg.org', 'lohrifestival.org', ['cultural and social history']]",23397776,"Require autoconfirmed or confirmed access (20:35, 4 August 2022)",136547,24 November 2001,Hagedis ,7109,18,2001-11-24,2001-11,2001
263,263,Estonia,https://en.wikipedia.org/wiki/Estonia,434,9,"['10.3176/arch.2012.supv1.11', '10.1787/9789264190801-en', '10.1093/biosci/bix014', '10.1007/978-94-6265-273-6', '10.2767/74735', '10.1038/s41467-020-19493-3', 'org/10.1515/9783110885996', '10.1007/978-3-642-29615-4_2', '10.4054/demres.2018.38.38', None, None, '28608869', None, None, '33293507', None, None, None, None, None, '5451287', None, None, '7723057', None, None, None]","[['estonian journal of archaeology'], [' energy policies beyond iea countries '], ['bioscience'], ['[[t.m.c. asser instituut'], ['publications office of the european union '], ['nature communications'], ['degruyter mouton '], ['[[springer publishing', (' lecture notes in computer science', ' science', 'science', 'v')], ['[[demographic research ']]",40,6,0,65,0,2,312,0.09216589861751152,0.013824884792626729,0.1497695852534562,0.020737327188940093,0.0,0.12672811059907835,9,"['finland.usembassy.gov', 'www.census.gov', 'dfat.gov', 'www.cia.gov', 'www.e-resident.gov', 'cia.gov', 'euobserver.com', 'www.estonianfreepress.com', 'books.google.com', 'www.google.com', 'www.nytimes.com', 'estonianworld.com', 'nordpoolspot.com', 'neweuropeaneconomy.com', 'books.google.com', 'www.newscientist.com', 'books.google.com', 'www.economist.com', 'books.google.com', 'www.alphr.com', 'books.google.com', 'www.prosperity.com', 'credit-suisse.com', 'www.reuters.com', 'www.gallup.com', 'qz.com', 'www.bbc.com', 'www.irishtimes.com', 'books.google.com', 'www.visitestonia.com', 'www.baltictimes.com', 'books.google.com', 'www.worldinfozone.com', 'www.yahoo.com', 'dw.com', 'mus-col.com', 'www.irishtimes.com', 'www.tasteatlas.com', 'estonianworld.com', 'lulu.com', 'www.wsj.com', 'www.wired.com', 'www.cnbc.com', 'www.worldinfozone.com', 'www.britannica.com', 'www.economist.com', 'www.bbc.com', 'books.google.com', 'www.google.com', 'balticbusinessnews.com', 'todellinentallinna.blogspot.com', 'books.google.com', 'www.bbc.com', 'kr-asia.com', 'www.economist.com', 'www.baltictimes.com', 'bachtrack.com', 'www.investinestonia.com', 'estonianworld.com', 'www.bbc.com', 'www.bbc.com', 'treasurytoday.com', 'estonianworld.com', '2020.stateofeuropeantech.com', 'www.gallup.com', 'books.google.com', 'www.country-studies.com', 'www.topuniversities.com', 'www.globalpolitician.com', 'e-estonia.com', 'www.cnbc.com', 'www.estonica.org', 'taxfoundation.org', 'www.oecd.org', 'www.doingbusiness.org', 'rsf.org', 'hdr.undp.org', 'data.worldbank.org', 'stats.oecd.org', 'www.norden.org', 'estonica.org', 'www.oecd.org', 'estonica.org', 'nordefco.org', 'lutheranworld.org', 'oikoumene.org', 'www.nordplusonline.org', 'www.oecd.org', 'www.oecd.org', 'www.fraserinstitute.org', 'www.estonica.org', 'www.pewforum.org', 'www.oecdbetterlifeindex.org', 'www.educationestonia.org', 'www.estonica.org', 'www.imf.org', 'assets.pewresearch.org', 'pewforum.org', 'www.world-nuclear-news.org', 'heritage.org', 'transparency.org', 'legacarta.intracen.org', 'www.nb8businessmobility.org', 'www.e3g.org', 'en.rsf.org', 'www.nrdc.org', 'www.wto.org', 'traceminternational.org', 'www.osce.org', 'www.osce.org', 'hdr.undp.org', ['estonian journal of archaeology'], [' energy policies beyond iea countries '], ['bioscience'], ['[[t.m.c. asser instituut'], ['publications office of the european union '], ['nature communications'], ['degruyter mouton '], ['[[springer publishing', (' lecture notes in computer science', ' science', 'science', 'v')], ['[[demographic research ']]",28222445,Require administrator access (no expiry set),239277,12 November 2001,134.132.88.xxx ,10405,23,2001-11-12,2001-11,2001
264,264,Mangaloreans,https://en.wikipedia.org/wiki/Mangaloreans,16,0,[],[],0,0,0,10,0,0,6,0.0,0.0,0.625,0.0,0.0,0.0,0,"['2fwww.daijiworld.com', 'www.hindu.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.daijiworld.com', 'www.hindu.com', 'info:q1h0nsiwwiej:scholar.google.com', 'www.hindu.com', 'www.newindianexpress.com', 'info:ytwrhamusnij:scholar.google.com']",20660037,Allow all users (no expiry set),21045,12 December 2008,Kensplanet ,468,3,2008-12-12,2008-12,2008
265,265,Kannur,https://en.wikipedia.org/wiki/Kannur,69,0,[],[],6,11,0,28,0,0,24,0.08695652173913043,0.15942028985507245,0.4057971014492754,0.0,0.0,0.2463768115942029,0,"['kannur.keralapolice.gov', 'lsgkerala.gov', 'imdpune.gov', 'mahe.gov', 'censusindia.gov', 'imdpune.gov', 'trend.kerala.gov', 'kannur.keralapolice.gov', 'censusindia.gov', 'kannurcorporation.lsgkerala.gov', 'censusindia.gov', 'www.timesnownews.com', 'indiarailinfo.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'www.facebook.com', 'www.thehindu.com', 'books.google.com', 'www.arabnews.com', 'books.google.com', 'books.google.com', 'deccanchronicle.com', 'ananthapuri.com', 'www.thehindu.com', 'www.bbc.com', 'www.facesplacesandplates.com', 'www.thehindu.com', 'economictimes.indiatimes.com', 'books.google.com', 'calicutnet.com', 'books.google.com', 'www.thehindu.com', 'www.thetakeiteasychef.com', 'www.deccanherald.com', 'www.thehindu.com', 'www.thehindu.com', 'www.timesnownews.com', 'indiarailinfo.com', 'www.cartage.org', 'urbanaffairskerala.org', 'www.keralatourism.org', 'www.kudumbashree.org', 'urbanaffairskerala.org', 'urbanaffairskerala.org']",2340298,Require administrator access (no expiry set),54777,30 July 2005,Nichalp ,2467,3,2005-07-30,2005-07,2005
266,266,Devon,https://en.wikipedia.org/wiki/Devon,89,0,[],[],7,16,0,11,0,0,55,0.07865168539325842,0.1797752808988764,0.12359550561797752,0.0,0.0,0.25842696629213485,0,"['www.devon.gov', 'www.ons.gov', 'www.northdevon.gov', 'www.gov', 'www.devon.gov', 'www.neighbourhood.statistics.gov', 'www.devon.gov', 'devon.gov', 'www.plymouth.gov', 'www.exmoor-nationalpark.gov', 'www.ons.gov', 'devon.gov', 'www.devon.gov', 'www.devon.gov', 'www.devon.gov', 'www.devon.gov', 'www.britannica.com', 'books.google.com', 'www.britannica.com', 'britannia.com', 'www.nature.com', 'www.christianitytoday.com', 'www.christianitytoday.com', 'www.gwr.com', 'variety.com', 'www.oxforddnb.com', 'users.senet.com', 'naturalengland.org', 'species.nbnatlas.org', 'www.devonbirds.org', 'www.northumbriacommunity.org', 'species.nbnatlas.org', 'plymouth-diocese.org', 'designatedsites.naturalengland.org']",8166,Require administrator access (no expiry set),83482,8 October 2001,212.248.133.xxx ,3095,6,2001-10-08,2001-10,2001
267,267,Islam in Kerala,https://en.wikipedia.org/wiki/Islam_in_Kerala,87,10,"['10.2307/2800388', '10.33306/mjssh/31', '10.5040/9780755610259.ch-013', '10.4324/9781003084129-11', '10.1159/000153449', '10.1017/9789048501069.008', '10.1163/22879811-12340009', None, None, None, None, '6745953', None, None, None, None, None, None, None, None, None]","[['man', 'royal anthropological institute of great britain and ireland'], ['muallim journal of social sciences and humanities'], ['i.b.tauris'], ['routledge'], ['human heredity'], ['global indian diasporas'], ['asian review of world histories']]",4,1,0,39,0,0,33,0.04597701149425287,0.011494252873563218,0.4482758620689655,0.11494252873563218,0.0,0.1724137931034483,7,"['censusindia.gov', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.frontlineonnet.com', 'www.thehindu.com', 'www.youtube.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'www.youtube.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'www.cookawesome.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thetakeiteasychef.com', 'books.google.com', 'www.facesplacesandplates.com', 'books.google.com', 'www.frontlineonnet.com', 'www.outlookindia.com', 'books.google.com', 'books.google.com', 'www.hindu.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.kozhikodeairport.com', 'books.google.com', 'worldcat.org', 'www.alislam.org', 'www.gutenberg.org', 'worldcat.org', ['man', 'royal anthropological institute of great britain and ireland'], ['muallim journal of social sciences and humanities'], ['i.b.tauris'], ['routledge'], ['human heredity'], ['global indian diasporas'], ['asian review of world histories']]",6172999,Allow all users (no expiry set),52697,29 July 2006,Shijaz ,510,0,2006-07-29,2006-07,2006
268,268,Saudi Arabia,https://en.wikipedia.org/wiki/Saudi_Arabia,688,10,"['10.1017/s0020743800028750', '10.1080/01436597.2021.1948325', '10.1186/s40985-019-0112-4', '10.1155/2012/642187', '10.1111/0020-8833.00053', '10.1038/s41598-021-89489-6', '10.1093/biosci/bix014', '10.1111/gwao.12626', '10.1038/news.2011.55', '10.1126/science.1199113', None, None, '30858991', '22523673', None, '33980918', '28608869', None, None, '21273486', None, None, '6391748', '3317126', None, '8115331', '5451287', None, None, None]","[['international journal of middle east studies '], ['third world quarterly'], ['public health reviews'], ['journal of nutrition and metabolism'], ['[[international studies quarterly'], ['scientific reports'], ['bioscience'], ['gender'], ['nature'], ['science ', 'science news ']]",91,41,0,256,0,32,259,0.13226744186046513,0.059593023255813955,0.37209302325581395,0.014534883720930232,0.0,0.2063953488372093,10,"['www.mofa.gov', 'www.state.gov', 'stats.gov', 'stats.gov', 'cia.gov', 'data.bls.gov', 'stats.gov', 'www.uscirf.gov', 'www.cia.gov', 'eia.doe.gov', 'www.cia.gov', 'stats.gov', 'laws.boe.gov', 'www.loc.gov', 'www.state.gov', '2009-2017.state.gov', '2001-2009.state.gov', 'www.moe.gov', 'stats.gov', 'stats.gov', 'stats.gov', 'www.state.gov', 'www.state.gov', 'eia.gov', 'www.eia.doe.gov', 'www.cia.gov', 'www.cia.gov', 'memory.loc.gov', '2009-2017.state.gov', '2001-2009.state.gov', 'www.state.gov', 'cia.gov', 'cia.gov', 'www.moe.gov', '2009-2017.state.gov', 'stats.gov', 'www.state.gov', 'stats.gov', 'www.cia.gov', 'www.mofa.gov', 'stats.gov', 'www.economist.com', 'www.wsj.com', 'www.economist.com', 'twitter.com', 'www.arabnews.com', 'www.ft.com', 'paleolithic-neolithic.com', 'www.reuters.com', 'chronicle.com', 'www.arabnews.com', 'books.google.com', 'www.arabnews.com', 'www.economist.com', 'www.thenationalnews.com', 'www.washingtonpost.com', 'www.smh.com', 'www.businessweek.com', 'www.bbc.com', 'arabnews.com', 'www.bbc.com', 'books.google.com', 'twitter.com', 'amp.cnn.com', 'www.nytimes.com', 'mirrorherald.com', 'www.nybooks.com', 'www.washingtonpost.com', 'www.cnbc.com', 'www.nationalgeographic.com', 'greenprophet.com', 'al-bab.com', 'arabianbusiness.com', 'www.economist.com', 'www.youtube.com', 'www.investopedia.com', 'www.reuters.com', 'www.cbsnews.com', 'www.nationthailand.com', 'saudigazette.com', 'uk.reuters.com', 'www.arabnews.com', 'books.google.com', 'ireport.cnn.com', 'selwaalhazzaa.com', 'news.nationalgeographic.com', 'variety.com', 'www.aljazeera.com', 'www.salon.com', 'twitter.com', 'www.economist.com', 'deadline.com', 'www.bloomberg.com', 'news.nationalgeographic.com', 'www.washingtonpost.com', 'books.google.com', 'www.washingtonpost.com', 'latimesblogs.latimes.com', 'www.thedailybeast.com', 'www.arabnews.com', 'www.thenationalnews.com', 'www.bbc.com', 'www.slate.com', 'www.saudiarabiatourismguide.com', 'www.thehindu.com', 'www.nytimes.com', 'www.elopak.com', 'www.bloomberg.com', 'todor66.com', 'books.google.com', 'america.aljazeera.com', 'www.arabnews.com', 'insidesaudi.com', 'www.arabnews.com', 'www.metrocorpcounsel.com', 'www.economist.com', 'www.businessinsider.com', 'www.bloomberg.com', 'arabnews.com', 'www.nybooks.com', 'country-stats.com', 'www.economist.com', 'www.voanews.com', 'bloomberg.com', 'www.time.com', 'www.economist.com', 'www.nbcnews.com', 'uk.reuters.com', 'books.google.com', 'www.montrealgazette.com', 'articles.cnn.com', 'www.britannica.com', 'archive.aramcoworld.com', 'www.nytimes.com', 'www.ipsos.com', 'www.ft.com', 'www.usatoday.com', 'www.al-monitor.com', 'www.britannica.com', 'www.nybooks.com', 'www.aljazeera.com', 'www.nytimes.com', 'news.vice.com', 'www.ft.com', 'www.hiiraan.com', 'www.economist.com', 'asiatimes.com', 'www.youtube.com', 'stepfeed.com', 'www.nytimes.com', 'www.christianpost.com', 'www.middleeastmonitor.com', 'books.google.com', 'mirrorherald.com', 'economictimes.indiatimes.com', 'www.atimes.com', 'books.google.com', 'www.newsweek.com', 'www.washingtonpost.com', 'www.albawaba.com', 'gulfnews.com', 'www.aljazeera.com', 'books.google.com', 'observers.france24.com', 'www.theglobeandmail.com', 'www.reuters.com', 'books.google.com', 'www.saudigazette.com', 'www.arabnews.com', 'books.google.com', 'www.nytimes.com', 'www.maritime-executive.com', 'www.bloomberg.com', 'ameinfo.com', 'deadline.com', 'www.businessinsider.com', 'www.washingtonpost.com', 'www.salon.com', 'books.google.com', 'arabnews.com', 'books.google.com', 'www.economist.com', 'www.reuters.com', 'thediplomat.com', 'pages.eiu.com', 'www.washingtonpost.com', 'arabnews.com', 'edition.cnn.com', 'www.arabnews.com', 'www.saudigazette.com', 'arabnews.com', 'www.saudigazette.com', 'news.yahoo.com', 'www.bloomberg.com', 'www.nytimes.com', 'www.youtube.com', 'www.time.com', 'www.washingtonpost.com', 'res.mdpi.com', 'www.nytimes.com', 'arabnews.com', 'www.theatlantic.com', 'res.mdpi.com', 'www.nytimes.com', 'www.wsj.com', 'www.reuters.com', 'www.reuters.com', 'www.nytimes.com', 'www.britannica.com', 'www.thepeninsulaqatar.com', 'www.arabnews.com', 'www.world-grain.com', 'www.aljazeera.com', 'www.nytimes.com', 'www.youtube.com', 'www.politico.com', 'books.google.com', 'www.arabnews.com', 'economist.com', 'books.google.com', 'books.google.com', 'arabianbusiness.com', 'www.economist.com', 'www.arabnews.com', 'books.google.com', 'www.saudigazette.com', 'abcnews.go.com', '2fwww.washingtonpost.com', 'www.natureindex.com', 'nostatusquo.com', 'aawsat.com', 'www.huffingtonpost.com', 'alriyadh.com', 'www.uidergisi.com', 'mondovisione.com', 'www.vice.com', 'www.economist.com', 'www.bbc.com', 'www.arabnews.com', 'arabianbusiness.com', 'www.bbc.com', 'www.dw.com', 'www.shanghairanking.com', 'cnn.com', 'books.google.com', 'www.mcclatchydc.com', 'www.businessinsider.com', 'ukessays.com', 'books.google.com', 'www.dailystar.com', 'www.newstatesman.com', 'www.washingtonpost.com', 'nasdaq.com', 'www.bloomberg.com', 'www.ethnologue.com', 'bloomberg.com', 'peakoil.com', 'books.google.com', 'books.google.com', 'www.economist.com', 'books.google.com', 'topics.nytimes.com', 'www.arabnews.com', 'docs.cdn.yougov.com', 'www.bloomberg.com', 'www.reuters.com', 'www.cnn.com', 'www.arabnews.com', 'www.cnbc.com', 'www.defensenews.com', 'www.reuters.com', 'arabnews.com', 'tdctrade.com', 'books.google.com', 'gulfnews.com', 'www.latimes.com', 'www.arriyadh.com', 'www.bbc.com', 'usatoday.com', 'www.britannica.com', 'www.reuters.com', 'www.economist.com', 'almodarresi.com', 'books.google.com', 'www.nytimes.com', 'www.middleeastmonitor.com', 'books.google.com', 'books.google.com', 'books.google.com', 'lebanonspring.com', 'time.com', 'foreignpolicy.com', 'www.wsj.com', 'www.economist.com', 'www.washingtonpost.com', 'www.bloomberg.com', 'www.nytimes.com', 'www.sipri.org', 'www.washingtoninstitute.org', 'arabstates.undp.org', 'worldfocus.org', 'whc.unesco.org', 'hdr.undp.org', 'www.cato.org', 'esa.un.org', 'weekly.ahram.org', 'memri.org', 'www.newsecuritybeat.org', 'www.sipri.org', 'www.pewforum.org', 'fas.org', 'persecutionofahmadis.org', 'whc.unesco.org', 'www.opec.org', 'www.us-sabc.org', 'nationalgeographic.org', 'www.meforum.org', 'whc.unesco.org', 'en.unesco.org', 'www.freedomhouse.org', 'www.wes.org', 'www.wssinfo.org', 'ich.unesco.org', 'pewforum.org', 'data.worldbank.org', 'data.worldbank.org', 'www.catsg.org', 'www.fishbase.org', 'www.un.org', 'www.catsg.org', 'www.transparency.org', 'opec.org', 'data.worldbank.org', 'sacm.org', 'globalsecurity.org', 'whc.unesco.org', 'www.npr.org', 'www.revealnews.org', 'www.freedomhouse.org', 'fas.org', 'jcpa.org', 'uis.unesco.org', 'www.unhcr.org', 'www.iiss.org', 'www.imf.org', 'carnegieendowment.org', 'www.globalsecurity.org', 'freedomhouse.org', 'memri.org', 'assets.pewresearch.org', 'www.jcpa.org', 'www.hrw.org', 'www.secularism.org', 'www.sipri.org', 'www.hrw.org', 'www.pbs.org', 'washwatch.org', 'www.un.org', 'hosted.ap.org', 'weekly.ahram.org', 'www.iags.org', 'npr.org', 'unstats.un.org', 'www.pewforum.org', 'whc.unesco.org', 'www.muhammadanism.org', 'data.worldbank.org', 'freedomhouse.org', 'sacm.org', 'sipri.org', 'www.pewforum.org', 'www.hrw.org', 'freedomhouse.org', 'www.amnesty.org', 'www.pewforum.org', 'www.amnesty.org', 'www.islamicpluralism.org', 'www.sciencemag.org', 'www.yemenileopard.org', 'www.pbs.org', 'www.cfr.org', 'hdr.undp.org', 'whc.unesco.org', 'www.newsecuritybeat.org', 'www.hrw.org', 'www.hrw.org', 'www.jstor.org', 'whc.unesco.org', ['international journal of middle east studies '], ['third world quarterly'], ['public health reviews'], ['journal of nutrition and metabolism'], ['[[international studies quarterly'], ['scientific reports'], ['bioscience'], ['gender'], ['nature'], ['science ', 'science news ']]",349303,Require autoconfirmed or confirmed access (no expiry set),327782,27 May 2001,KoyaanisQatsi ,13033,24,2001-05-27,2001-05,2001
269,269,Province of Avellino,https://en.wikipedia.org/wiki/Province_of_Avellino,3,0,[],[],0,0,0,0,0,0,3,0.0,0.0,0.0,0.0,0.0,0.0,0,[],1418064,Allow all users (no expiry set),7219,21 January 2005,Markussep ,195,0,2005-01-21,2005-01,2005
270,270,Republic of Ireland,https://en.wikipedia.org/wiki/Republic_of_Ireland,296,4,"['10.1093/obo/9780199846719-0149', '10.1093/biosci/bix014', '10.1086/424697', '10.1086/508399', None, '28608869', '15309688', None, None, '5451287', '1182057', None]","[[' oxford university press '], ['bioscience'], ['am. j. hum. genet. '], ['journal of british studies']]",22,8,0,78,0,3,182,0.07432432432432433,0.02702702702702703,0.2635135135135135,0.013513513513513514,0.0,0.11486486486486487,4,"['www.cia.gov', 'www.budget.gov', 'www.agriculture.gov', 'www.taoiseach.gov', 'www.cia.gov', 'taoiseach.gov', 'www.cia.gov', 'www.inis.gov', 'books.google.com', '2fwww.irishtimes.com', 'www.irishtimes.com', 'books.google.com', 'www.bloomberg.com', 'www.irishtimes.com', 'www.irishtimes.com', '2fwww.irishtimes.com', 'irishcentral.com', 'www.irishtimes.com', 'www.afl.com', 'www.irishtimes.com', '247wallst.com', 'www.irishtimes.com', 'www.latimes.com', 'books.google.com', 'cbonds.com', '2fwww.irishtimes.com', 'www.irishtimes.com', 'www.irishexaminer.com', 'www.irishtimes.com', 'www1.skysports.com', 'turnerscross.com', 'www.ft.com', 'books.google.com', 'wesleyjohnston.com', 'www.irishtimes.com', 'www.megalithomania.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.irishtimes.com', 'travelinireland.com', 'www.reuters.com', 'www.irelandlogue.com', 'www.irishtimes.com', 'www.ulsterscotsagency.com', 'www.forbes.com', 'www.irishtimes.com', 'books.google.com', 'www.irishtimes.com', 'www.irishexaminer.com', '2fwww.irishtimes.com', 'books.google.com', 'www.irishtimes.com', 'www.worldgolf.com', 'www.irishtimes.com', 'www.irishtimes.com', 'www.irishtimes.com', 'www.rugbyleagueplanet.com', 'www.idaireland.com', 'nationmaster.com', 'www.historyireland.com', 'www.bloomberg.com', '2fonline.wsj.com', 'www.irishtimes.com', 'www.healthpowerhouse.com', 'crwflags.com', 'www.irishtimes.com', 'books.google.com', 'www.irishtimes.com', 'www.irishtimes.com', 'books.google.com', 'www.irishtimes.com', 'books.google.com', 'about.com', 'www.irishtimes.com', 'books.google.com', 'www.idaireland.com', 'newsfeed.time.com', 'www.latimes.com', 'www.bbc.com', 'ballybegvillage.com', 'www.ft.com', 'www.cbsnews.com', 'www.finance-magazine.com', '2fwww.irishtimes.com', 'www.irishtimes.com', 'oecdbetterlifeindex.org', 'worldtimelines.org', 'www.nyulawglobal.org', 'worldtimelines.org', 'www.secularism.org', 'www.worldlii.org', 'www.secularism.org', 'hdr.undp.org', 'hdr.undp.org', 'www.imf.org', 'www.catholicculture.org', 'imf.org', 'www.worldcat.org', 'hbr.org', 'www.oecd.org', 'www.iata.org', 'treaties.un.org', 'www.nyulawglobal.org', 'www.catholicculture.org', 'oecd.org', 'ourworldindata.org', 'www.ancientfortresses.org', [' oxford university press '], ['bioscience'], ['am. j. hum. genet. '], ['journal of british studies']]",14560,Require administrator access (no expiry set),228280,14 October 2001,213.122.201.xxx ,11894,21,2001-10-14,2001-10,2001
271,271,San Marino,https://en.wikipedia.org/wiki/San_Marino,83,2,"['10.1093/biosci/bix014', '10.1038/s41467-020-19493-3', '28608869', '33293507', '5451287', '7723057']","[['bioscience'], ['nature communications']]",11,3,0,33,0,1,33,0.13253012048192772,0.03614457831325301,0.39759036144578314,0.024096385542168676,0.0,0.1927710843373494,2,"['www.gov', 'www.cia.gov', 'history.state.gov', 'www.lonelyplanet.com', 'books.google.com', 'www.sanmarinosite.com', 'www.nytimes.com', 'www.everyculture.com', 'sanmarinosite.com', 'scoreshelf.com', 'm.youtube.com', 'www.mister-baseball.com', 'www.publibook.com', 'www.reuters.com', 'espnfc.com', 'www.washingtonpost.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.bbc.com', 'www.sanmarinosite.com', 'www.visitsanmarino.com', 'sanmarinosite.com', 'sanmarinosite.com', 'sanmarinosite.com', 'newsweek.com', 'weatherspark.com', 'books.google.com', 'politifact.com', 'rtwin30days.com', 'www.visitsanmarino.com', 'www.thoughtco.com', 'int.soccerway.com', 'jewishencyclopedia.com', 'sports.yahoo.com', 'www.venditafrancobolli.com', 'ais-sanmarino.org', 'imf.org', 'www.fao.org', 'imf.org', 'www.bandamilitaresanmarino.org', 'www.unescap.org', 'newadvent.org', 'jewishvirtuallibrary.org', 'www.unece.org', 'climate-data.org', 'pubdocs.worldbank.org', ['bioscience'], ['nature communications']]",27248,Require autoconfirmed or confirmed access (no expiry set),78444,27 May 2001,KoyaanisQatsi ,3886,19,2001-05-27,2001-05,2001
272,272,Kenya,https://en.wikipedia.org/wiki/Kenya,272,12,"['10.1017/s0022278x00016657', '10.1017/s0022278x00000082', '10.1080/02604027.2014.894868', '10.1017/s0022278x00003980', '10.1080/17531055.2020.1863642', '10.1126/science.aao2646', '10.2307/220649', '10.2307/1160687', '10.1093/afraf/adg007', '10.1038/s41467-020-19493-3', '10.1353/at.1999.0008', '10.1353/arw.2012.0010', None, None, None, None, None, '29545508', None, None, None, '33293507', None, None, None, None, None, None, None, None, None, None, None, '7723057', None, None]","[[' the journal of modern african studies '], ['the journal of modern african studies'], ['world futures'], [' the journal of modern african studies'], ['journal of eastern african studies'], ['science'], ['the international journal of african historical studies'], [' africa'], [' african affairs '], ['nature communications'], ['africa today'], ['african studies review']]",54,9,0,62,0,5,130,0.19852941176470587,0.03308823529411765,0.22794117647058823,0.04411764705882353,0.0,0.2757352941176471,12,"['2001-2009.state.gov', 'www.usaid.gov', 'www.cia.gov', 'cia.gov', 'www.parliament.vic.gov', 'www.loc.gov', 'lcweb2.loc.gov', '2009-2017.state.gov', 'www.cia.gov', 'www.constructionkenya.com', 'www.quakerinfo.com', 'businessdailyafrica.com', 'www.chimpreports.com', 'ngm.nationalgeographic.com', 'nationsencyclopedia.com', 'www.nytimes.com', 'www.supersport.com', 'www.businessdailyafrica.com', 'www.businessdailyafrica.com', 'www.britannica.com', 'en-maktoob.news.yahoo.com', 'www.time.com', 'ethnologue.com', 'www.kenyatraveltips.com', 'www.thoughtco.com', 'www.bbc.com', 'howwemadeitinafrica.com', 'www.bbc.com', 'www.nytimes.com', 'swahilihub.com', 'www.theautochannel.com', 'www.ft.com', 'www.ft.com', 'kapsowarhospital.com', 'worldnews.nbcnews.com', 'dhsprogram.com', 'magicalkenya.com', 'www.highbeam.com', 'empowermentopportunities.com', 'indcatholicnews.com', 'af.reuters.com', 'www.aljazeera.com', 'www.nytimes.com', 'www.yellowpageskenya.com', 'africanews.com', 'www.kenyaembassy.com', 'www.reuters.com', 'www.bbc.com', 'www.nytimes.com', 'www.climatestotravel.com', 'www.theatlantic.com', 'www.railjournal.com', 'www.businessdailyafrica.com', 'www.business-anti-corruption.com', 'www.nytimes.com', 'www.washingtonpost.com', 'www.bloomberg.com', 'www.bloomberg.com', 'www.washingtonpost.com', 'www.csmonitor.com', 'news.nationalgeographic.com', 'af.reuters.com', 'www.google.com', 'www.cnn.com', 'www.reuters.com', 'archive.fiba.com', 'www.chimpreports.com', 'edition.cnn.com', 'www.africanews.com', 'www.bbc.com', 'orvillejenkins.com', 'archive.ipu.org', 'www.unaids.org', 'data.worldbank.org', 'www.climatelinks.org', 'transparency.org', 'www.npr.org', 'www.ediec.org', 'kenyaconstitution.org', 'www.irinnews.org', 'hdr.undp.org', 'www.pbs.org', 'unhcr.org', 'kenyaun.org', 'pewglobal.org', 'www.pbs.org', 'data.worldbank.org', 'imf.org', 'worldbank.org', 'www.norrag.org', 'www.worldbank.org', 'www.knchr.org', 'www.mfi-upgrading-initiative.org', 'exploreit.icrisat.org', 'www.ilo.org', 'unicef.org', 'kenyalaw.org', 'www.imf.org', 'www.unhcr.org', 'nationalgeographic.org', 'www.wfp.org', 'data.worldbank.org', 'www.womenconnect.org', 'www.cipe.org', 'phdtree.org', 'www.pewglobal.org', 'imf.org', 'www.iea.org', 'www.britishmuseum.org', 'www.amnesty.org', 'wrfnet.org', 'imf.org', 'www.kenyalaw.org', 'cdkn.org', 'conferences.ifpri.org', 'racism.org', 'kenya.opendataforafrica.org', 'kenyaconnection.org', 'www.pbs.org', 'unstats.un.org', 'oikoumene.org', 'www.doingbusiness.org', 'globalsecurity.org', 'www.pbs.org', 'unstats.un.org', [' the journal of modern african studies '], ['the journal of modern african studies'], ['world futures'], [' the journal of modern african studies'], ['journal of eastern african studies'], ['science'], ['the international journal of african historical studies'], [' africa'], [' african affairs '], ['nature communications'], ['africa today'], ['african studies review']]",188171,Require administrator access (no expiry set),203512,1 November 2001,208.60.199.xxx ,9332,16,2001-11-01,2001-11,2001
273,273,Uttarakhand,https://en.wikipedia.org/wiki/Uttarakhand,134,1,"['10.1007/s13659-019-0202-5', '30968350', '6538708']",[['natural products and bioprospecting']],16,13,0,62,0,0,42,0.11940298507462686,0.09701492537313433,0.4626865671641791,0.007462686567164179,0.0,0.22388059701492538,1,"['www.censusindia.gov', 'censusindia.gov', 'schooleducation.uk.gov', 'censusindia.gov', 'transport.uk.gov', 'schooleducation.uk.gov', 'www.censusindia.gov', 'censusindia.gov', 'planningcommission.gov', 'uk.gov', 'nfdb.gov', 'censusindia.gov', 'schooleducation.uk.gov', 'www.whatismyresults.com', 'www.business-standard.com', 'euttaranchal.com', 'www.ndtv.com', 'www.gmvnl.com', 'twitter.com', 'www.india-today.com', 'uttaraguide.com', 'www.telegraphindia.com', 'bedupako.com', 'zeenews.india.com', 'www.collinsdictionary.com', 'www.jagran.com', 'www.thehindu.com', 'www.lonelyplanet.com', 'articles.timesofindia.indiatimes.com', 'www.indianexpress.com', 'corbett-national-park.com', 'm.timesofindia.com', 'humaribaat.com', 'indianexpress.com', 'www.ethnologue.com', 'www.voatibetanenglish.com', 'books.google.com', 'www.jagranjosh.com', 'books.google.com', 'www.jagran.com', 'timesofindia.indiatimes.com', 'm.economictimes.com', 'www.outlookindia.com', 'www.dailypioneer.com', 'books.google.com', 'www.business-standard.com', 'www.tribuneindia.com', 'www.hindustantimes.com', 'www.jankarihub.com', 'www.britannica.com', 'articles.timesofindia.indiatimes.com', 'statisticstimes.com', 'aboututtarakhand.com', 'www.livehindustan.com', 'www.quora.com', 'www.jagran.com', 'books.google.com', 'www.euttarakhand.com', 'books.google.com', 'pppinindia.com', 'lonelyplanet.com', 'timesofindia.indiatimes.com', 'www.tribuneindia.com', 'www.timesnownews.com', 'www.mapsofindia.com', 'dictionary.reference.com', 'uttaranchal-india.com', 'www.collinsdictionary.com', 'www.tribuneindia.com', 'www.thehindu.com', 'www.hindustantimes.com', 'www.nainitaltourism.com', 'www.lonelyplanet.com', 'www.amarujala.com', 'www.hindustantimes.com', 'www.unesco.org', 'hdr.undp.org', 'whc.unesco.org', 'whc.unesco.org', 'ich.unesco.org', 'www.ibef.org', 'uttarakhandforest.org', 'www.devalsari.org', 'www.iisd.org', 'www.unesco.org', 'hdi.globaldatalab.org', 'www.downtoearth.org', 'www.unesco.org', 'www.downtoearth.org', 'impactfactor.org', 'www.unesco.org', ['natural products and bioprospecting']]",1429154,Allow all users (no expiry set),116313,25 January 2005,Ceti ,5178,27,2005-01-25,2005-01,2005
274,274,Odisha,https://en.wikipedia.org/wiki/Odisha,144,1,"['10.1038/nindia.2019.69', None, None]",[['nature india ']],10,23,0,86,0,0,24,0.06944444444444445,0.1597222222222222,0.5972222222222222,0.006944444444444444,0.0,0.2361111111111111,1,"['lawodisha.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'censusindia.gov', 'odisha.gov', 'nfdb.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'www.odisha.gov', 'www.wildlife.odisha.gov', 'www.archive.india.gov', 'odishapolice.gov', 'www.odisha.gov', 'magazines.odisha.gov', 'www.imd.gov', 'www.orissa.gov', 'www.censusindia.gov', 'odisha.gov', 'www.censusindia.gov', 'stscodisha.gov', 'www.censusindia.gov', 'odisha.gov', 'magazines.odisha.gov', 'www.pragativadi.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.telegraphindia.com', 'books.google.com', 'www.thehindubusinessline.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'www.telegraphindia.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.dnaindia.com', 'kalingatv.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'www.newindianexpress.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.orissalinks.com', 'books.google.com', 'news.webindia123.com', 'www.goal.com', 'www.newindianexpress.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.newindianexpress.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'www.ndtv.com', 'books.google.com', 'www.simplytadka.com', 'books.google.com', 'www.thehindu.com', 'www.dailypioneer.com', 'books.google.com', 'timesofindia.indiatimes.com', 'odissi.itgo.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'indianexpress.com', 'ibnlive.in.com', 'www.newindianexpress.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'www.dailypioneer.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.jagranjosh.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'www.financialexpress.com', 'rediff.com', 'www.dailypioneer.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.rediff.com', 'books.google.com', 'www.prsindia.org', 'www.unesco.org', 'globaldatalab.org', 'www.assocham.org', 'hdi.globaldatalab.org', 'globaldatalab.org', 'www.worldbank.org', 'www.seaturtle.org', 'www.bput.org', 'www.wwfindia.org', ['nature india ']]",250724,Require administrator access (no expiry set),126735,21 June 2003,Cyberagent ,6890,4,2003-06-21,2003-06,2003
275,275,Balearic Islands,https://en.wikipedia.org/wiki/Balearic_Islands,56,4,"['10.1093/zoolinnean/zlaa094', '10.1016/j.quaint.2007.06.039', '10.1038/s41559-020-1102-0', '10.1007/s10963-008-9010-2', None, None, '32094539', None, None, None, '7080320', None]","[['zoological journal of the linnean society'], ['quaternary international'], ['nature ecology '], ['journal of world prehistory']]",2,0,0,12,0,0,38,0.03571428571428571,0.0,0.21428571428571427,0.07142857142857142,0.0,0.10714285714285714,4,"['www.vice.com', 'directferries.com', 'www.magentayachts.com', 'rsssf.com', 'www.magentayachts.com', 'books.google.com', 'rsssf.com', 'www.lavanguardia.com', 'majorcadailybulletin.com', 'www.andalucia-for-holidays.com', 'www.hellenicaworld.com', 'sobreespana.com', 'www.eoearth.org', 'www.mantleplumes.org', ['zoological journal of the linnean society'], ['quaternary international'], ['nature ecology '], ['journal of world prehistory']]",21336521,Require administrator access (no expiry set),53324,20 May 2002,Jeronimo ,1456,3,2002-05-20,2002-05,2002
276,276,Slovenia,https://en.wikipedia.org/wiki/Slovenia,339,5,"['10.1177/0959683610371998', '10.1038/s41467-020-19493-3', '10.1093/biosci/bix014', '10.1007/s10531-012-0246-x', '10.7152/ssj.v12i1.3797', None, '33293507', '28608869', None, None, None, '7723057', '5451287', None, None]","[['the holocene '], ['nature communications'], ['bioscience'], [' biodiversity and conservation '], [' slovene studies journal']]",21,28,0,60,0,1,224,0.061946902654867256,0.08259587020648967,0.17699115044247787,0.014749262536873156,0.0,0.1592920353982301,5,"['mo.gov', 'www.arso.gov', 'www.cia.gov', 'www.gov', 'natura2000.gov', 'ukom.gov', 'www.cia.gov', 'kazalci.arso.gov', 'www.ukom.gov', 'www.svz.gov', 'www.arso.gov', 'mop.gov', 'mop.gov', 'www.arso.gov', 'arso.gov', 'kazalci.arso.gov', 'mzp.gov', 'www.zgs.gov', 'mop.gov', 'www.cia.gov', 'www.zgs.gov', 'ukom.gov', '.gov', 'www.arso.gov', 'www.ukom.gov', 'www.mss.gov', 'kazalci.arso.gov', 'arhiv.mm.gov', 'books.google.com', 'www.sloveniatimes.com', 'books.google.com', 'www.collinsdictionary.com', 'books.google.com', 'www.economist.com', 'www.geodetski-vestnik.com', 'olympiandatabase.com', 'www.nationalgeographic.com', 'www.geodetski-vestnik.com', 'www.bbc.com', 'books.google.com', 'worldcasinodirectory.com', 'www.britannica.com', 'ngm.nationalgeographic.com', 'balkan-trout.com', 'books.google.com', 'books.google.com', 'www.cnbc.com', 'www.kozina.com', 'books.google.com', 'mladinska.com', 'books.google.com', 'books.google.com', 'docs.google.com', 'sloveniatimes.com', 'www.theslovenian.com', 'www.nogomania.com', 'books.google.com', 'www.sloveniatimes.com', 'seenews.com', 'www.shanghairanking.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.sloveniatimes.com', 'books.google.com', 'earthinpictures.com', 'books.google.com', 'www.sloveniatimes.com', 'books.google.com', 'www.bloomberg.com', 'books.google.com', 'vecer.com', 'books.google.com', 'www.britannica.com', 'www.infoplease.com', 'www.everyculture.com', 'books.google.com', 'books.google.com', 'books.google.com', 'arising-empire.com', 'webcache.googleusercontent.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'www.total-slovenia-news.com', 'books.google.com', 'www.sloveniatimes.com', 'books.google.com', 'oecdbetterlifeindex.org', 'www.porttechnology.org', 'europeanregionofgastronomy.org', 'data.worldbank.org', 'www.oecd.org', 'documents.worldbank.org', 'whc.unesco.org', 'www.morigenos.org', 'imf.org', 'data.oecd.org', 'communistcrimes.org', 'www.heritage.org', 'imf.org', 'www.oecd.org', 'communistcrimes.org', 'zacat.gesis.org', 'www.wilsoncenter.org', 'jewishvirtuallibrary.org', 'hdr.undp.org', 'www.olympic.org', 'www.fao.org', ['the holocene '], ['nature communications'], ['bioscience'], [' biodiversity and conservation '], [' slovene studies journal']]",27338,Require administrator access (no expiry set),235770,27 May 2001,KoyaanisQatsi ,9274,22,2001-05-27,2001-05,2001
277,277,Ancient Egypt,https://en.wikipedia.org/wiki/Ancient_Egypt,116,10,"['10.1038/ncomms15694', '10.1136/bmj.e8268', None, '10.1111/j.1469-1809.2008.00493.x', '10.2307/1356573', '10.2307/3822337', '10.1002/ajpa.20569', '10.1016/j.jasrep.2017.12.025', '10.3390/genes9030135', '10.1086/371778', '28556824', '23247979', '23888738', '19053990', None, None, '17295300', None, '29494531', None, '5459999', None, None, None, None, None, None, None, '5867856', None]","[[' nature communications '], ['bmj'], ['medicinski pregled'], [' annals of human genetics '], ['[[bulletin of the american schools of oriental research'], ['[[journal of egyptian archaeology'], ['[[american journal of physical anthropology'], [' journal of archaeological science'], ['genes'], ['[[journal of near eastern studies']]",8,0,0,53,0,1,44,0.06896551724137931,0.0,0.45689655172413796,0.08620689655172414,0.0,0.15517241379310345,10,"['books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.livescience.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.nbcnews.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'edition.cnn.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'discovermagazine.com', 'books.google.com', 'books.google.com', 'seeker.com', 'books.google.com', 'archive.archaeology.org', 'www.eoearth.org', 'www.metmuseum.org', 'www.archaeology.org', 'www.britishmuseum.org', 'www.reshafim.org', 'www.worldcat.org', 'mysteriousuniverse.org', [' nature communications '], ['bmj'], ['medicinski pregled'], [' annals of human genetics '], ['[[bulletin of the american schools of oriental research'], ['[[journal of egyptian archaeology'], ['[[american journal of physical anthropology'], [' journal of archaeological science'], ['genes'], ['[[journal of near eastern studies']]",874,Require administrator access (no expiry set),138970,13 May 2001,LA2 ,7998,2,2001-05-13,2001-05,2001
278,278,Armenians,https://en.wikipedia.org/wiki/Armenians,120,7,"['10.1038/ejhg.2011.192', '10.1017/s0010417520000432', '10.5281/zenodo.1240524', '10.1038/ejhg.2015.206', '10.11606/issn.2763-650x.i6p109-115', '10.1515/if-2018-0009', '22085901', None, None, '26486470', None, None, '3286660', None, None, '4820045', None, None]","[[' european journal of human genetics '], ['comparative studies in society and history'], [''], ['european journal of human genetics'], ['revista de estudos orientais'], ['indogermanische forschungen', 'the university of british columbia library']]",6,5,0,25,0,0,77,0.05,0.041666666666666664,0.20833333333333334,0.058333333333333334,0.0,0.15,6,"['diaspora.gov', 'mniejszosci.narodowe.mac.gov', 'www.immi.gov', 'www.ukrcensus.gov', 'www.stat.gov', 'www.tacentral.com', 'armenianweekly.com', 'oglobo.globo.com', 'books.google.com', 'books.google.com', 'www.todayszaman.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.armdiasporamuseum.com', 'armenianow.com', 'books.google.com', 'www.reuters.com', 'books.google.com', 'www.britannica.com', 'www.nytimes.com', 'books.google.com', 'www.tacentral.com', 'www.worldinfozone.com', 'www.ncccusa.org', 'www.holyland.org', 'www.armenialiberty.org', 'www.anca.org', 'sino-platonic.org', 'www.armenialiberty.org', [' european journal of human genetics '], ['comparative studies in society and history'], [''], ['european journal of human genetics'], ['revista de estudos orientais'], ['indogermanische forschungen', 'the university of british columbia library']]",387816,Require autoconfirmed or confirmed access (no expiry set),91226,4 December 2003,145.254.191.241 ,4396,13,2003-12-04,2003-12,2003
279,279,Lithuanians,https://en.wikipedia.org/wiki/Lithuanians,48,5,"['10.1371/journal.pone.0135820', '10.1016/j.cub.2019.04.026', '10.1001/archpedi.158.1.27', '10.1086/320123', '26332464', '31080083', '14706954', '11309683', '4558026', '6544527', None, '1226098', 'ncbi']","[['plos one '], ['current biology '], [' archives of pediatrics '], [' [[the american journal of human genetics'], 'ncbi']",1,6,0,7,0,0,29,0.020833333333333332,0.125,0.14583333333333334,0.10416666666666667,0.0,0.25,5,"['osp.stat.gov', 'db1.stat.gov', 'osp.stat.gov', 'factfinder.census.gov', 'www.stat.gov', 'www.dhs.gov', 'epoca.globo.com', 'www.britannica.com', 'de.statista.com', 'www.khazaria.com', 'ltuworld.com', 'www.britannica.com', 'www.ltuworld.com', 'lituanus.org', ['plos one '], ['current biology '], [' archives of pediatrics '], [' [[the american journal of human genetics'], 'ncbi']",459375,Allow all users (no expiry set),44804,7 February 2004,Altenmann ,1521,15,2004-02-07,2004-02,2004
280,280,Tamil Nadu,https://en.wikipedia.org/wiki/Tamil_Nadu,271,4,"['10.1353/asi.2003.0031', '10.1017/s0021911807001234', '10.2307/2943246', '10.2307/2053325', None, None, None, None, None, None, None, None]","[['asian perspectives '], ['the journal of asian studies '], ['the journal of asian studies '], ['the journal of asian studies ']]",20,32,0,129,0,1,85,0.07380073800738007,0.11808118081180811,0.47601476014760147,0.014760147601476014,0.0,0.2066420664206642,4,"['www.tnpolice.gov', 'www.tn.gov', 'ennoreport.gov', 'censusindia.gov', 'mnre.gov', 'censusindia.gov', 'www.tn.gov', 'ddindia.gov', 'www.tourism.gov', 'www.tnrd.gov', 'www.tn.gov', 'censusindia.gov', 'www.censusindia.gov', 'www.tn.gov', 'www.tnpolice.gov', 'indcom.tn.gov', 'india.gov', 'www.censusindia.gov', 'cbfcindia.gov', 'www.tn.gov', 'www.tnrd.gov', 'tourism.gov', 'censusindia.gov', 'www.tn.gov', 'assembly.tn.gov', 'www.censusindia.gov', 'tn.gov', 'www.tn.gov', 'www.tn.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'pibmumbai.gov', 'www.hindu.com', 'economictimes.indiatimes.com', 'tamilnadu.com', 'www.thehindu.com', 'www.thenewsminute.com', 'books.google.com', 'www.thehindu.com', 'britannica.com', 'www.aishtma.com', 'www.openthemagazine.com', 'www.thenewsminute.com', 'www.thehindubusinessline.com', 'www.espncricinfo.com', 'www.thehindu.com', 'books.google.com', 'www.crayondata.com', 'www.thehindu.com', 'www.newindianexpress.com', 'articles.timesofindia.indiatimes.com', 'books.google.com', 'www.espncricinfo.com', 'books.google.com', 'rediff.com', 'www.thehindu.com', 'www.hinduonnet.com', 'theswaddle.com', 'www.hinduonnet.com', 'books.google.com', 'www.nytimes.com', 'articles.timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'winentrance.com', 'www.financialexpress.com', 'www.thehindubusinessline.com', 'www.thehindu.com', 'news.google.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.business-standard.com', 'books.google.com', 'www.hindu.com', 'www.historynet.com', 'www.thenewsminute.com', 'www.espncricinfo.com', 'www.espncricinfo.com', 'museumstuff.com', 'timesofindia.indiatimes.com', 'media.daimler.com', 'www.hindu.com', 'mapsofindia.com', 'www.winentrance.com', 'www.indiantelevision.com', 'outlookindia.com', 'www.britannica.com', 'www.espncricinfo.com', 'www.rediff.com', 'www.thehindu.com', 'www.washingtonpost.com', 'aljazeera.com', 'www.espncricinfo.com', 'archive.financialexpress.com', 'www.hindu.com', 'www.hindu.com', 'yamaha-motor-india.com', 'www.newindianexpress.com', 'economictimes.indiatimes.com', 'shadowchief.com', 'www.newslaundry.com', 'www.shanlax.com', 'www.espncricinfo.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'www.newindianexpress.com', 'www.hindu.com', 'www.thehindu.com', 'books.google.com', 'www.resourceinvestor.com', 'timesofindia.indiatimes.com', 'www.hindu.com', 'www.jio.com', 'www.hindu.com', 'blessingsonthenet.com', 'prabinsamuel.medium.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'indianexpress.com', 'www.hindu.com', 'www.thehindu.com', 'www.hindu.com', 'articles.timesofindia.indiatimes.com', 'www.deccanchronicle.com', 'www.findcollegereviews.com', 'www.financialexpress.com', 'timesofindia.indiatimes.com', 'www.hindu.com', 'timesofindia.indiatimes.com', 'www.hindu.com', 'www.hindu.com', 'www.tndte.com', 'www.thehindu.com', 'www.openthemagazine.com', 'tamilnadu.com', 'books.google.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'www.dnaindia.com', 'www.thehindu.com', 'teauction.com', 'www.thehindu.com', 'books.google.com', 'www.thehindubusinessline.com', 'tamilnadu.com', 'www.thehindu.com', 'articles.timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'tamilnadu.com', 'www.eximfile.com', 'articles.timesofindia.indiatimes.com', 'www.hathway.com', 'articles.timesofindia.indiatimes.com', 'www.uniindia.com', 'www.thehindu.com', 'www.hindu.com', 'www.ibef.org', 'globaldatalab.org', 'www.ibef.org', 'whc.unesco.org', 'www.ciil-classicaltamil.org', 'unesdoc.unesco.org', 'hdrstats.undp.org', 'tnhighways.org', 'whc.unesco.org', 'www.rubberboard.org', 'mssrf.org', 'whc.unesco.org', 'www.hindunet.org', 'tamilculturewaterloo.org', 'unsystem.org', 'siteresources.worldbank.org', 'asc-india.org', 'www.sciencenews.org', 'assets.wwfindia.org', 'www.sriaurobindoashram.org', ['asian perspectives '], ['the journal of asian studies '], ['the journal of asian studies '], ['the journal of asian studies ']]",29918,Require extended confirmed access (no expiry set),189323,18 August 2001,24.108.233.xxx ,12604,7,2001-08-18,2001-08,2001
281,281,Malta,https://en.wikipedia.org/wiki/Malta,334,16,"['10.1017/s0003598x00097787', '10.3406/camed.1998.1231', '10.2307/296290', '10.1023/a:1005386004103', '10.1093/biosci/bix014', 'gov.mt/en/islands/dates.asp', '10.2307/621508', 'gov.mt', '10.1080/09518960412331302203', '10.1016/j.cities.2004.07.001', '10.3233/jrs-1996-9104', '10.1136/jramc-138-03-09', '10.5281/zenodo.1181783', '10.1023/a:1006888926016', '10.3390/resources7030058', None, None, None, None, '28608869', None, None, None, None, None, '23512022', '1453384', None, None, None, None, None, None, None, '5451287', None, None, None, None, None, None, None, None, None, None]","[['antiquity '], ['cahiers de la méditerranée '], ['journal of roman studies '], ['international journal for the advancement of counselling'], ['bioscience '], ['department of information'], ['transactions of the institute of british geographers '], ['doi.gov.mt'], ['mediterranean historical review '], ['cities '], ['international journal of risk '], ['journal of the royal army medical corps '], ['language science press '], ['geojournal '], ['resources ']]",33,38,0,140,0,1,106,0.09880239520958084,0.11377245508982035,0.41916167664670656,0.04790419161676647,0.0,0.26047904191616766,15,"['nso.gov', 'privatisation.gov', 'sahha.gov', 'docs.justice.gov', 'mitc.gov', 'www.nso.gov', 'www.creativemalta.gov', 'www.gov', 'nso.gov', '2001-2009.state.gov', 'afm.gov', 'nso.gov', 'www.nso.gov', 'privatisation.gov', 'www.cia.gov', 'www.gov', 'justiceservices.gov', 'www.gov', 'dossier.ogp.noaa.gov', 'www.gov', 'nso.gov', 'www.metoffice.gov', 'privatisation.gov', 'afm.gov', 'afm.gov', 'agriculture.gov', 'www.lc.gov', 'privatisation.gov', 'www.cia.gov', 'foreignaffairs.gov', 'www.cia.gov', 'www.royal.gov', 'justiceservices.gov', 'www.culturalheritage.gov', 'www.nso.gov', 'nso.gov', 'www.nso.gov', 'nso.gov', 'www.euractiv.com', 'www.tns-opinion.com', 'www.maltatoday.com', 'www.geocities.com', 'timesofmalta.com', 'encarta.msn.com', 'www.cnn.com', 'www.dailymalta.com', 'apartments.com', 'silentrebellion.newsvine.com', 'www.britannica.com', 'books.google.com', 'www.timesofmalta.com', 'www.bbc.com', 'www.tvm.com', 'www.pressreader.com', 'www.maltairport.com', 'www.independent.com', 'www.timesofmalta.com', 'melitensiawth.com', 'timesofmalta.com', 'www.timesofmalta.com', 'www.independent.com', 'weatherbase.com', 'aboutmalta.com', 'books.google.com', 'www.timesofmalta.com', 'visitmalta.com', 'www.libyaherald.com', 'books.google.com', 'books.google.com', 'maltaramc.com', 'www.supernovamalta.com', 'www.timesofmalta.com', 'books.google.com', 'www.timesofmalta.com', 'books.google.com', 'books.google.com', 'www.biblegateway.com', 'www.independent.com', 'www.maltastreetmap.com', 'books.google.com', 'aapa.files.cms-plus.com', 'timesofmalta.com', 'archive.maltatoday.com', 'www.independent.com', 'www.independent.com', 'timesofmalta.com', 'books.google.com', 'maltatoday.com', 'books.google.com', 'www.aboutmalta.com', 'books.google.com', 'www.timesofmalta.com', 'www.bloomberg.com', 'books.google.com', 'www.timesofmalta.com', 'www.trofeocaza.com', 'www.independent.com', 'www.timesofmalta.com', 'www.maltadata.com', 'www.trofeocaza.com', 'www.independent.com', 'www.timesofmalta.com', 'www.petroleumafrica.com', 'hopeandoptimism.com', 'www.napoleonicsociety.com', 'maltaweathersite.com', 'books.google.com', 'books.google.com', 'www.timesofmalta.com', 'melitensiawth.com', 'www.malta.com', 'books.google.com', 'www.dw.com', 'www.timesofmalta.com', 'www.timesofmalta.com', 'books.google.com', 'alloexpat.com', 'www.timesofmalta.com', 'www.timesofmalta.com', 'www.timesofmalta.com', 'www.independent.com', 'www.timesofmalta.com', 'books.google.com', 'www.maltavoyager.com', 'bay.com', 'www.gozoandmalta.com', 'books.google.com', 'indexmundi.com', 'environmentalgraffiti.com', 'books.google.com', 'archive.maltatoday.com', 'www.weather2travel.com', 'www.melitensiawth.com', 'www.maltawildplants.com', 'www.nationmaster.com', 'maltaweather.com', 'articles.latimes.com', 'www.clevelandjewishnews.com', 'visitmalta.com', 'edrichton.com', 'www.visitmalta.com', 'www.timesofmalta.com', 'www.airmalta.com', 'encyclopedia2.thefreedictionary.com', 'www.maltatoday.com', 'buddeblog.com', 'www.maltamigration.com', 'macmillandictionaries.com', 'books.google.com', 'www.independent.com', 'visitmalta.com', 'www.pressreader.com', 'elpais.com', 'www.britannica.com', 'lulu.com', 'www.timesofmalta.com', 'knoema.com', 'jimdiamondmd.com', 'www.independent.com', 'www.aboutmalta.com', 'geocities.com', 'icef.com', 'books.google.com', 'tripadvisor.com', 'www.maltaculture.com', 'maltaweather.com', 'www.independent.com', 'timesofindia.indiatimes.com', 'newsbook.com', 'books.google.com', 'www.visitmalta.com', 'maltatoday.com', 'carnaval.com', 'www.di-ve.com', 'www.malta-tix.com', 'www.maltauncovered.com', 'www.timesofmalta.com', 'www.independent.com', 'www.newadvent.org', 'data.footprintnetwork.org', 'whc.unesco.org', 'www.scubed.org', 'www.pvv.org', 'financemalta.org', 'www.hrw.org', 'www.financemalta.org', 'www.un.org', 'www.imf.org', 'www.localhistories.org', 'otsf.org', 'treaties.un.org', 'unwto.org', 'seatemperature.org', 'imf.org', 'www.inta-aivn.org', 'culturemalta.org', 'www.patrimonju.org', 'centralbankmalta.org', 'otsf.org', 'www.centralbankmalta.org', 'www.micc.org', 'www.islandofgozo.org', 'whc.unesco.org', 'ictsamalta.org', 'www.stbenedictcollege.org', 'www.mca.org', 'hdr.undp.org', 'meteo-climat-bzh.dyndns.org', 'era.org', 'whc.unesco.org', 'gerom.org', ['antiquity '], ['cahiers de la méditerranée '], ['journal of roman studies '], ['international journal for the advancement of counselling'], ['bioscience '], ['department of information'], ['transactions of the institute of british geographers '], ['doi.gov.mt'], ['mediterranean historical review '], ['cities '], ['international journal of risk '], ['journal of the royal army medical corps '], ['language science press '], ['geojournal '], ['resources ']]",19137,Require administrator access (no expiry set),246395,20 May 2001,KoyaanisQatsi ,11045,47,2001-05-20,2001-05,2001
282,282,North Indian culture,https://en.wikipedia.org/wiki/North_Indian_culture,3,0,[],[],1,0,0,1,0,0,1,0.3333333333333333,0.0,0.3333333333333333,0.0,0.0,0.3333333333333333,0,"['www.culturenorthindia.com', 'whc.unesco.org']",32866391,Allow all users (no expiry set),13217,25 August 2011,Greatbuddha ,261,2,2011-08-25,2011-08,2011
283,283,Hangzhou,https://en.wikipedia.org/wiki/Hangzhou,122,4,"['10.1787/9789264230040-en', '10.1163/9789004366152_008', '10.1126/science.1166605', '10.1017/s0041977x02000320', None, None, '19299619', None, None, None, None, None]","[['[[organisation for economic co-operation and development'], ['brill '], [' science '], ['bulletin of the school of oriental and african studies']]",7,10,0,52,0,0,49,0.05737704918032787,0.08196721311475409,0.4262295081967213,0.03278688524590164,0.0,0.1721311475409836,4,"['www.zj.gov', 'zjjcmspublic.oss-cn-hangzhou-zwynet-d01-a.internet.cloud.zj.gov', 'hzindus.gov', 'old-cdc.cma.gov', 'museum.shqp.gov', 'www.zj.stats.gov', 'www.hangzhou.gov', 'hmc.hz.gov', 'cdc.cma.gov', 'www.ehangzhou.gov', 'china-window.com', 'www.timeshighereducation.com', 'www.topuniversities.com', 'www.theborneopost.com', 'www.yhwt.com', 'books.google.com', 'time.com', 'www.washingtonpost.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.ssdph.com', 'hangzhou.com', 'jewish-holiday.com', 'www.usnews.com', 'www.docin.com', 'www.demographia.com', 'hangzhouweekly.com', 'www.schiphol.com', 'www.dailyexpress.com', 'books.google.com', 'www.natureindex.com', 'www.minorsights.com', 'www.shanghairanking.com', 'www.docin.com', 'www.scmp.com', 'chinaautoweb.com', 'www.fjnet.com', 'www.joneslanglasalle.com', 'www.chinatoday.com', 'books.google.com', 'news.xinhuanet.com', 'bbs.hangzhou.com', 'www.natureindex.com', 'www.china-briefing.com', 'ori.hangzhou.com', 'www.time.com', 'www.channelnewsasia.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.pwccn.com', 'news.sina.com', 'www.tellerreport.com', 'geography.about.com', 'www.nbcnews.com', 'www.chinapages.com', 'www.zj.xinhuanet.com', 'time.com', 'hangzhou.zjol.com', 'news.xinhuanet.com', 'www.un.org', 'www.china.org', 'china.org', 'www.mherrera.org', 'kotakinabalu.china-consulate.org', 'www.chinaheritagequarterly.org', 'www.china.org', ['[[organisation for economic co-operation and development'], ['brill '], [' science '], ['bulletin of the school of oriental and african studies']]",158185,Allow all users (no expiry set),111047,15 December 2002,Roadrunner ,2570,5,2002-12-15,2002-12,2002
284,284,Lithuania,https://en.wikipedia.org/wiki/Lithuania,502,8,"['10.1038/s41467-020-19493-3', '10.1046/j.1529-8817.2003.00119.x', '10.5194/hess-7-423-2003', '10.1038/s41467-018-02825-9', '10.1057/palgrave.fp.8200087', '10.1093/biosci/bix014', '10.1038/d41586-018-05308-5', '33293507', '15469421', None, '29382937', None, '28608869', '29872189', '7723057', None, None, '5789860', None, '5451287', None]","[['nature communications'], ['annals of human genetics '], ['hydrology and earth system sciences '], ['nature communications'], ['french politics ', '[[palgrave macmillan'], ['bioscience'], ['nature']]",60,17,0,68,0,1,348,0.11952191235059761,0.03386454183266932,0.13545816733067728,0.01593625498007968,0.0,0.1693227091633466,7,"['osp.stat.gov', 'state.gov', 'www.cia.gov', 'www.cia.gov', 'osp.stat.gov', 'www.cia.gov', 'www.cia.gov', 'osp.stat.gov', 'www.cia.gov', 'www.osac.gov', 'osp.stat.gov', 'osp.stat.gov', 'state.gov', 'osp.stat.gov', 'osp.stat.gov', 'ops.stat.gov', 'www.stat.gov', 'statista.com', 'euractiv.com', 'www.statista.com', 'books.google.com', 'baltictimes.com', 'sites.google.com', 'www.youtube.com', 'travel-earth.com', 'investlithuania.com', 'books.google.com', 'fdiintelligence.com', 'www.bloomberg.com', 'www.ft.com', 'www.britannica.com', 'www.wired.com', 'www.bloomberg.com', 'www.credit-suisse.com', 'www.vanlifetribe.com', 'books.google.com', 'books.google.com', 'nasdaqbaltic.com', 'enterpriselithuania.com', 'voanews.com', 'www.eshopworld.com', 'books.google.com', 'www.britannica.com', 'whiteguide-nordic.com', 'wtvbam.com', 'books.google.com', 'urbanadventures.com', 'media.daimler.com', 'www.bbc.com', 'books.google.com', 'truelithuania.com', 'geosite.jankrogh.com', 'maistologija.wordpress.com', 'books.google.com', 'www.nytimes.com', 'public.dhe.ibm.com', 'uptimeinstitute.com', 'books.google.com', 'books.google.com', 'books.google.com', 'investlithuania.com', 'hoophall.com', 'baltic-course.com', 'pr.nba.com', 'www.youtube.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'wtvbam.com', 'flandersinvestmentandtrade.com', 'lonelyplanet.com', 'www.volvogroup.com', 'www.euronews.com', 'books.google.com', 'thebalance.com', 'lightcon.com', 'www.bbc.com', 'www.foreignaffairs.com', 'books.google.com', 'cloudscene.com', 'fatbirder.com', 'books.google.com', 'www.fdiintelligence.com', 'global.truelithuania.com', 'crowdfundinsider.com', 'oecd.org', 'www.yadvashem.org', 'www.european-agency.org', 'lituanus.org', 'wayback.archive-it.org', 'www.oecd.org', 'childmortality.org', 'whc.unesco.org', 'www.imf.org', 'lituanus.org', 'www.bdforum.org', 'wttc.org', 'unesdoc.unesco.org', 'data.worldbank.org', 'gpseducation.oecd.org', 'www.imf.org', 'data.oecd.org', 'publicadministration.un.org', 'publicadministration.un.org', 'brewersofeurope.org', 'lituanus.org', 'partizanai.org', 'www.ushmm.org', 'ich.unesco.org', 'partizanai.org', 'data.oecd.org', 'theeuropeanlibrary.org', 'umc.org', 'www.lituanus.org', 'data.oecd.org', 'www.partizanai.org', 'www.wto.org', 'web.arcive.org', 'stats.oecd.org', 'oecd.org', 'www.imf.org', 'devdata.worldbank.org', 'm.epo.org', 'childmortality.org', 'www.constituteproject.org', 'lituanus.org', 'www.imf.org', 'www3.weforum.org', 'un.org', 'draugas.org', 'www.partizanai.org', 'datahelpdesk.worldbank.org', 'unstats.un.org', 'www.draugas.org', 'climate-change-performance-index.org', 'healthmanagement.org', 'w3.unece.org', 'www.partizanai.org', 'hdr.undp.org', 'world-nuclear.org', 'wits.worldbank.org', 'www.currency-iso.org', 'bellona.org', 'partizanai.org', 'lokashakti.org', ['nature communications'], ['annals of human genetics '], ['hydrology and earth system sciences '], ['nature communications'], ['french politics ', '[[palgrave macmillan'], ['bioscience'], ['nature']]",17675,Require administrator access (no expiry set),307381,17 April 2001,BruceMiller ,11245,32,2001-04-17,2001-04,2001
285,285,Luxembourg,https://en.wikipedia.org/wiki/Luxembourg,236,2,"['10.1093/acrefore/9780190228637.013.1041', '10.1038/s41467-020-19493-3', None, '33293507', None, '7723057']","[['oxford university press'], ['nature communications']]",17,9,0,30,0,2,176,0.07203389830508475,0.038135593220338986,0.1271186440677966,0.00847457627118644,0.0,0.11864406779661017,2,"['www.treasury.gov', 'www.cia.gov', 'www.cia.gov', 'www.sepb.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.treasury.gov', 'www.cia.gov', 'www.com', 'www.railjournal.com', 'www.telx.com', 'www.henleypassportindex.com', 'www.sprooch.com', 'escxtra.com', 'www.britannica.com', 'pwc.com', 'www.ft.com', 'www.economist.com', 'www.telx.com', 'soluxions-magazine.com', 'stadiumdb.com', 'netindex.com', 'shenandoahdavis.canalblog.com', 'www.britannica.com', 'www.britannica.com', 'www.worldatlas.com', 'www.atlasandboots.com', 'www.hollywoodreporter.com', 'www.eiu.com', 'www.britannica.com', 'financialsecrecyindex.com', 'tns-ilres.com', 'countryeconomy.com', 'www.bloomberg.com', 'www.fidomes.com', 'www.britannica.com', 'www.britannica.com', 'uptimeinstitute.com', 'www.imf.org', 'www.migrationinformation.org', 'www.nizkor.org', 'www.oecd.org', 'imf.org', 'www.globalinnovationindex.org', 'healthmanagement.org', 'whc.unesco.org', 'zacat.gesis.org', 'whc.unesco.org', 'hdr.undp.org', 'www.un.org', 'stats.oecd.org', 'www.heritage.org', 'features.pewforum.org', 'globalsecurity.org', 'stats.oecd.org', ['oxford university press'], ['nature communications']]",17515,Require administrator access (no expiry set),134496,17 May 2001,Pinkunicorn ,6349,12,2001-05-17,2001-05,2001
286,286,Assyrian people,https://en.wikipedia.org/wiki/Assyrian_people,339,18,"['10.1086/373570', '10.3378/1534-6617(2008)80[73:vodvaa]2.0.co;2', '10.1111/j.1354-5078.2000.00363.x', '10.1086/511103', None, '10.1086/677249', '10.22425/jul.2004.5.1.1', '10.1371/journal.pone.0187408', '10.3109/03014460.2010.535562', '10.1093/hgs/dcz045', '10.1163/157338406780345899', '10.1371/journal.pone.0041252', '10.7227/bjrl.78.3.14', '10.1163/22118993-90000037', '10.2307/1797632', '10.1038/81685', None, None, None, None, '3456196', None, None, '29099847', '21329477', None, None, '22815981', None, None, None, '11062480', None, None, None, None, '1684716', None, None, '5669434', None, None, None, '3399854', None, None, None, None]","[['journal of near eastern studies'], ['hum biol '], [' [[nations and nationalism '], ['journal of near eastern studies'], [' american journal of human genetics '], ['journal of near eastern studies'], ['journal of universal language'], ['plos one'], ['ann. hum. biol. '], ['holocaust and genocide studies'], ['iran and the caucasus '], [' plos one'], ['the bulletin of the john rylands library'], [' muqarnas'], ['the journal of the royal geographical society of london'], [' nature genetics ']]",57,9,0,144,0,0,111,0.168141592920354,0.02654867256637168,0.4247787610619469,0.05309734513274336,0.0,0.24778761061946902,16,"['factfinder.census.gov', 'factfinder2.census.gov', 'www.abs.gov', 'www.azleg.gov', 'www.state.gov', '2001.ukrcensus.gov', 'archive.stats.gov', 'www.state.gov', 'factfinder.census.gov', 'books.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'chaldeanflag.com', 'books.google.com', 'books.google.com', 'www.warscapes.com', 'books.google.com', 'books.google.com', 'www.hurriyetdailynews.com', 'www.syriacstudies.com', 'books.google.com', 'roadsandkingdoms.com', 'adherents.com', 'www.reuters.com', 'www.syriacsnews.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.christiansofiraq.com', 'books.google.com', 'crwflags.com', 'books.google.com', 'www.biomedcentral.com', 'books.google.com', 'www.trtworld.com', 'books.google.com', 'warscapes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.sbs.com', 'books.google.com', 'books.google.com', 'www.christianpost.com', 'www.trtworld.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'paloaltoonline.com', 'books.google.com', 'books.google.com', 'www.dailytelegraph.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.ethnologue.com', 'books.google.com', 'books.google.com', 'www.seyfocenter.com', 'www.astanatimes.com', 'dictionary.com', 'books.google.com', 'www.britannica.com', 'www.boston.com', 'books.google.com', 'britannica.com', 'books.google.com', 'armenianweekly.com', 'books.google.com', 'en.hawarnews.com', 'books.google.com', 'adherents.com', 'www.ishtartv.com', 'www.haaretz.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.al-monitor.com', 'warisboring.com', 'books.google.com', 'www.jokopost.com', 'diepresse.com', 'books.google.com', 'www.christianpost.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.france24.com', 'catholicphilly.com', 'books.google.com', 'www.al-monitor.com', 'www.fredaprim.com', 'www.qenshrin.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.usnews.com', 'www.nationalreview.com', 'www.jokopost.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'www.christianheadlines.com', 'books.google.com', 'www.atour.com', 'crwflags.com', 'books.google.com', 'www.al-monitor.com', 'parstimes.com', 'books.google.com', 'books.google.com', 'trackbill.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.todayszaman.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'syrianobserver.com', 'books.google.com', 'www.sbs.com', 'books.google.com', 'books.google.com', 'www.assyrianconference.com', 'gedsh.bethmardutho.org', 'zowaa.org', 'www.jaas.org', 'www.jaas.org', 'www.cpa-iraq.org', 'www.unhcr.org', 'www.aleteia.org', 'aina.org', 'peshitta.org', 'www.assyrianpolicy.org', 'www.aina.org', 'www.newadvent.org', 'aina.org', 'mag.jewishinseattle.org', 'aina.org', 'www.refworld.org', 'www.jaas.org', 'www.npr.org', 'www.jaas.org', 'www.aina.org', 'unpo.org', 'www.jaas.org', 'www.assyrianfoundation.org', 'www.ssi.org', 'syrianorthodoxchurch.org', 'www.jaas.org', 'en.wikisource.org', 'www.jstor.org', 'www.assyrianpolicy.org', 'www.jaas.org', 'www.jstor.org', 'www.nestorian.org', 'www.jaas.org', 'aina.org', 'aina.org', 'www.aina.org', 'www.assyrianpolicy.org', 'www.aina.org', 'www.culturalsurvival.org', 'www.iranicaonline.org', 'www.worldhistory.org', 'unpo.org', 'gedsh.bethmardutho.org', 'gedsh.bethmardutho.org', 'aanf.org', 'www.meforum.org', 'worldhistory.org', 'www.aina.org', 'www.aina.org', 'www.eurfedling.org', 'www.aina.org', 'www.assyrianpolicy.org', 'www.refworld.org', 'spectator.org', 'indict.org', 'www.aina.org', 'www.shlama.org', ['journal of near eastern studies'], ['hum biol '], [' [[nations and nationalism '], ['journal of near eastern studies'], [' american journal of human genetics '], ['journal of near eastern studies'], ['journal of universal language'], ['plos one'], ['ann. hum. biol. '], ['holocaust and genocide studies'], ['iran and the caucasus '], [' plos one'], ['the bulletin of the john rylands library'], [' muqarnas'], ['the journal of the royal geographical society of london'], [' nature genetics ']]",266350,Require administrator access (no expiry set),178543,13 July 2003,69.14.67.183 ,7659,8,2003-07-13,2003-07,2003
287,287,Castellabate,https://en.wikipedia.org/wiki/Castellabate,2,0,[],[],0,0,0,0,0,0,2,0.0,0.0,0.0,0.0,0.0,0.0,0,[],6125780,Allow all users (no expiry set),5439,26 July 2006,Dr. Blofeld ,119,0,2006-07-26,2006-07,2006
288,288,Berbers,https://en.wikipedia.org/wiki/Berbers,216,17,"['10.1086/386295', '10.1525/aa.1956.58.3.02a00390', '10.1080/13629380500409917', '10.1186/1471-2148-14-109', '10.1080/09503110.2019.1706372', '10.1371/journal.pgen.1004393.s017', '10.1093/jts/os-xliii.171-172.188', '10.1093/jss/xliii.2.209', '10.1126/science.306.5702.1680c', '10.1007/s00439-005-1266-3', '10.1086/386294', '10.1086/340669', '10.1086/423147', '10.1371/journal.pgen.1002397', '10.1073/pnas.1800851115', '10.1093/gbe/evv118', '15069642', None, None, '24885141', None, '24921250', None, None, '15576591', '15806398', '15042509', '11992266', '15202071', '22253600', '29895688', '26108492', '1181965', None, None, '4062890', None, '4055572', None, None, None, None, '1181964', '379148', '1216069', '3257290', '6042094', '4524485']","[['american journal of human genetics'], ['american anthropologist'], ['the journal of north african studies'], ['[[bmc evolutionary biology'], ['al-masāq'], ['[[plos genetics', 'plos genetics '], ['[[the journal of theological studies'], ['[[journal of semitic studies'], ['science'], ['human genetics'], ['american journal of human genetics'], ['american journal of human genetics'], ['american journal of human genetics'], ['[[plos genetics'], ['[[proceedings of the national academy of sciences'], ['[[genome biology and evolution']]",14,12,0,48,0,0,125,0.06481481481481481,0.05555555555555555,0.2222222222222222,0.0787037037037037,0.0,0.19907407407407407,16,"['www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'commune-mahdia.gov', 'www.census.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', '2001-2009.state.gov', 'www.cia.gov', 'www.cia.gov', '2001-2009.state.gov', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.google.com', 'books.google.com', 'books.google.com', 'www.christianitytoday.com', 'books.google.com', 'www.theglobeandmail.com', 'www.moroccoworldnews.com', 'www.foxnews.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'books.google.com', 'mondeberbere.com', 'news.vice.com', 'www.nytimes.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.wafin.com', 'books.google.com', 'www.aljazeera.com', 'www.elwatan.com', 'worldpopulationreview.com', 'www.aljazeera.com', 'www.washtimes.com', 'www.britannica.com', 'books.google.com', 'www.sfgate.com', 'lexicorient.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'sfgate.com', 'www.elwatan.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.langues-de-france.org', 'www.jstor.org', 'www.orthodoxengland.org', 'www.metmuseum.org', 'aaregistry.org', 'minorityrights.org', 'whc.unesco.org', 'en.wiktionary.org', 'www.newadvent.org', 'unpo.org', 'whc.unesco.org', 'journals.openedition.org', 'globalheritagefund.org', 'www.ccel.org', ['american journal of human genetics'], ['american anthropologist'], ['the journal of north african studies'], ['[[bmc evolutionary biology'], ['al-masāq'], ['[[plos genetics', 'plos genetics '], ['[[the journal of theological studies'], ['[[journal of semitic studies'], ['science'], ['human genetics'], ['american journal of human genetics'], ['american journal of human genetics'], ['american journal of human genetics'], ['[[plos genetics'], ['[[proceedings of the national academy of sciences'], ['[[genome biology and evolution']]",48132,Require administrator access (no expiry set),173735,7 April 2002,Pgdudda ,8303,16,2002-04-07,2002-04,2002
289,289,Serbs,https://en.wikipedia.org/wiki/Serbs,202,15,"['0350-0861/2014/0350-08611402099t.pdf', '10.2307/2498513', '10.2298/gei1301119s', '10.1016/j.gene.2012.01.030', '10.1371/journal.pone.0135820', '10.1163/19552629-01202003', '10.2298/eka1403029r', '10.1098/rsos.161054', '10.2298/pkjif1480203b', '10.1111/nana.12433', '10.1080/0963749022000009225', '10.1075/jlp.12.3.02ivk', '10.1080/00905990903239174', '10.1080/14690760600963198', None, None, None, '22310393', '26332464', None, None, '28484621', None, None, None, None, None, None, None, None, None, None, '4558026', None, None, '5414258', None, None, None, None, None, None]","[['glasnik etnografskog instituta sanu'], [' slavic review'], ['glasnik etnografskog instituta'], ['gene '], ['plos one '], ['journal of language contact '], ['economic annals'], ['royal society open science'], ['prilozi za knjizevnost i jezik'], [' journal of genocide research '], ['religion'], ['journal of language and politics', '[[john benjamins publishing company'], ['nationalities papers'], [' totalitarian movements and political religions']]",9,6,0,83,0,0,89,0.04455445544554455,0.0297029702970297,0.41089108910891087,0.07425742574257425,0.0,0.1485148514851485,14,"['factfinder2.census.gov', 'nasa.gov', 'www.siepa.gov', 'www.stat.gov', 'www.vti.mod.gov', 'www.immi.gov', 'books.google.com', 'scholar.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.atptour.com', 'books.google.com', 'books.google.com', 'www.ebritic.com', 'books.google.com', 'www.serbiaconsulatenyc.com', 'books.google.com', 'books.google.com', 'www.vreme.com', 'theculturetrip.com', 'books.google.com', 'www.atptour.com', 'books.google.com', 'www.idahostatesman.com', 'books.google.com', 'books.google.com', 'books.google.com', 'balkaninsight.com', 'books.google.com', 'www.nytimes.com', 'www.nba.com', 'books.google.com', 'mozzartsport.com', 'books.google.com', 'www.scribd.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'soccerlens.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.pregled-rs.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.scribd.com', 'books.google.com', 'books.google.com', 'www.nba.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.premierleague.com', 'www.merriamwebster.com', 'books.google.com', 'www.vreme.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'reuters.com', 'books.google.com', 'books.google.com', 'www.forbes.com', 'books.google.com', 'books.google.com', 'www.wtatennis.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.monstat.org', 'www.maticasrpska.org', 'www.unicef.org', 'royalfamily.org', 'www.yadvashem.org', 'www.eserbia.org', 'minorityrights.org', 'faostat.fao.org', 'www.monstat.org', ['glasnik etnografskog instituta sanu'], [' slavic review'], ['glasnik etnografskog instituta'], ['gene '], ['plos one '], ['journal of language contact '], ['economic annals'], ['royal society open science'], ['prilozi za knjizevnost i jezik'], [' journal of genocide research '], ['religion'], ['journal of language and politics', '[[john benjamins publishing company'], ['nationalities papers'], [' totalitarian movements and political religions']]",59512,Allow all users (no expiry set),124047,26 June 2002,Jeronimo ,6905,10,2002-06-26,2002-06,2002
290,290,Mango,https://en.wikipedia.org/wiki/Mango,85,26,"['10.5415/apallergy.2011.1.1.43', '10.3389/fpls.2017.00577', '10.1016/j.foodchem.2012.08.029', '10.1080/09637480410001666441', '10.1016/j.canlet.2008.01.047', '10.1016/j.plaphy.2010.02.012', '10.1016/j.foodchem.2008.09.107', '10.1111/j.0105-1873.2004.00451.x', '10.1038/sj.ejcn.1602841', '10.1016/j.foodchem.2011.06.053', '10.1021/jf800738r', '10.1007/978-94-011-1584-1_8', '10.1007/s11130-006-0035-3', '10.1111/j.0105-1873.2005.00454.x', '10.1016/s0021-9673(04)01406-2', '10.1016/j.abb.2005.05.015', None, '10.1016/j.phytochem.2010.05.024', '10.1111/nph.15731', '10.1016/j.plaphy.2013.07.006', '10.1136/bmj.297.6664.1639', '10.1186/s12870-015-0663-6', '10.1002/jsfa.3692', '10.1021/jf060566s', '10.1016/j.tplants.2020.01.005', '10.1021/jf0484069', '22053296', '28473837', '23122101', '14985189', '18359153', '20363641', None, '15606656', '17637601', None, '18558692', None, '17243011', '15701120', '15553152', '15979560', '11381849', '20598721', '30730057', '23911730', '3147776', '26573148', None, '16968105', '32191870', '15740041', '3206236', '5397511', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, '1838873', '4647706', None, None, None, None]","[['asia pacific allergy'], ['frontiers in plant science '], [' food chemistry'], ['int j food sci nutr '], ['cancer lett '], ['plant physiology and biochemistry'], [' food chemistry'], ['contact dermatitis '], ['eur j clin nutr '], [' food chemistry'], ['j agric food chem '], ['springer netherlands'], ['plant foods hum nutr '], ['contact dermatitis '], ['j chromatogr a '], ['arch biochem biophys '], ['cutis '], [' phytochemistry'], ['new phytologist '], [' plant physiology and biochemistry'], ['british medical journal '], ['bmc plant biology '], ['journal of the science of food and agriculture'], ['j agric food chem '], ['trends in plant science'], ['j agric food chem ']]",6,4,0,24,0,0,25,0.07058823529411765,0.047058823529411764,0.2823529411764706,0.3058823529411765,0.0,0.4235294117647059,26,"['india.gov', 'archive.india.gov', 'www.usaid.gov', 'www.usaid.gov', 'www.thestar.com', 'www.rappler.com', 'www.diariesofmagazine.com', 'rediff.com', 'www.thedailyrecords.com', 'travel.nytimes.com', 'www.marketmanila.com', 'www.telegraphindia.com', 'www.journalnow.com', 'www.exoticindiaart.com', 'toptropicals.com', 'bdnews24.com', 'www.arabnews.com', 'www.etymonline.com', 'in.lifestyle.yahoo.com', 'bdnews24.com', 'www.wheninmanila.com', 'www.springerplus.com', 'nmb-database.com', 'vahrehvah.com', 'www.sciencedirect.com', 'www.nytimes.com', 'www.thelittleepicurean.com', 'www.bdnews24.com', 'www.fao.org', 'www.crfg.org', 'www.fao.org', 'webexhibits.org', 'actahort.org', 'croplife.org', ['asia pacific allergy'], ['frontiers in plant science '], [' food chemistry'], ['int j food sci nutr '], ['cancer lett '], ['plant physiology and biochemistry'], [' food chemistry'], ['contact dermatitis '], ['eur j clin nutr '], [' food chemistry'], ['j agric food chem '], ['springer netherlands'], ['plant foods hum nutr '], ['contact dermatitis '], ['j chromatogr a '], ['arch biochem biophys '], ['cutis '], [' phytochemistry'], ['new phytologist '], [' plant physiology and biochemistry'], ['british medical journal '], ['bmc plant biology '], ['journal of the science of food and agriculture'], ['j agric food chem '], ['trends in plant science'], ['j agric food chem ']]",56315,Require administrator access (no expiry set),53178,12 June 2002,Stepnwolf ,8353,6,2002-06-12,2002-06,2002
291,291,Ancient Rome,https://en.wikipedia.org/wiki/Ancient_Rome,322,9,"['10.1086/367123', '10.1126/science.aay6826', '10.1086/367079', '10.1086/366973', '10.5195/jwsr.2006.369', '10.1126/science.366.6466.673', '10.2307/1170959', '10.1016/j.cub.2021.04.022', '10.1086/367078', None, '31699931', None, None, None, '31699914', None, '33974848', None, None, '7093155', None, None, None, None, None, None, None]","[['classical philology '], [' science'], ['classical philology '], ['classical philology'], ['journal of world-systems research'], ['[[science ', '[[american association for the advancement of science'], ['social science history'], ['current biology'], ['classical philology ']]",30,0,0,56,0,0,228,0.09316770186335403,0.0,0.17391304347826086,0.027950310559006212,0.0,0.12111801242236025,9,"['books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.bresciamusei.com', 'www.ancientlibrary.com', 'books.google.com', 'www.britannica.com', 'www.newyorker.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.bresciamusei.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.unrv.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'adriangoldsworthy.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'ancienthistory.about.com', 'www.britannica.com', 'books.google.com', 'www.amazon.com', 'books.google.com', 'warfarehistorynetwork.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.questia.com', 'books.google.com', 'www.huffingtonpost.com', 'books.google.com', 'books.google.com', 'www.highbeam.com', 'books.google.com', 'books.google.com', 'www.roman-emperors.org', 'www.roman-emperors.org', 'www.roman-emperors.org', 'www.historyguide.org', 'www.ibiblio.org', 'www.britishmuseum.org', 'www.gutenberg.org', 'www.gutenberg.org', 'www.worldhistory.org', 'www.gutenberg.org', 'www.metmuseum.org', 'www.historyguide.org', 'www.txclassics.org', 'www.roman-emperors.org', 'www.gutenberg.org', 'www.roman-emperors.org', 'livius.org', 'www.gutenberg.org', 'www.metmuseum.org', 'www.roman-emperors.org', 'library.thinkquest.org', 'www.roman-emperors.org', 'smarthistory.khanacademy.org', 'www.roman-emperors.org', 'www.roman-emperors.org', 'theottomans.org', 'www.roman-emperors.org', 'insidescience.org', 'www.gutenberg.org', 'livius.org', ['classical philology '], [' science'], ['classical philology '], ['classical philology'], ['journal of world-systems research'], ['[[science ', '[[american association for the advancement of science'], ['social science history'], ['current biology'], ['classical philology ']]",521555,Require administrator access (no expiry set),228398,12 March 2004,Muriel Gottrop~enwiki ,6429,12,2004-03-12,2004-03,2004
292,292,Lilium,https://en.wikipedia.org/wiki/Lilium,105,10,"['10.1270/jsbbs.52.207', '10.1016/j.ympev.2004.12.023', '10.1007/s00606-011-0524-1', '10.3389/fpls.2021.699226', '10.1016/0168-9452(91)90262-7', '10.2460/javma.2002.220.49', '10.1007/s00122-004-1739-0', '10.1270/jsbbs.51.39', '10.1053/j.tcam.2010.09.006', '10.1007/s00606-006-0513-y', None, '15878122', None, None, None, '12680447', '15290047', None, '21147474', None, None, None, None, None, None, None, None, None, None, None]","[['育種学雑誌 breeding science '], ['molecular phylogenetics and evolution'], ['plant systematics and evolution'], ['frontiers in plant science '], ['plant science '], ['j. am. vet. med. assoc. '], ['theoretical and applied genetics '], ['育種学雑誌 breeding science '], ['topics in companion animal medicine'], ['plant systematics and evolution ']]",20,10,0,32,0,0,33,0.19047619047619047,0.09523809523809523,0.3047619047619048,0.09523809523809523,0.0,0.38095238095238093,10,"['hdais.coa.gov', 'www.gov', 'consumer.fda.gov', 'www.mohw.gov', 'www.ops.gov', 'www.nbnky.gov', 'hdais.coa.gov', 'hdais.coa.gov', 'www.ops.gov', 'www.moh.gov', 'books.google.com', 'books.google.com', 'books.google.com', 'www.sohu.com', 'www.gardeners.com', 'books.google.com', 'homeguides.sfgate.com', 'www.perennials.com', 'www.teleflora.com', 'books.google.com', 'cpfd.cnki.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.perennials.com', 'www.vethelpdirect.com', 'www.libertytimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'brentandbeckysbulbs.com', 'www.buzzle.com', 'designresearchgroup.wordpress.com', 'www.elnuevodia.com', 'www.lemonlilyfestival.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.sunstar.com', 'www.aspcapro.org', 'efloras.org', 'efloras.org', 'lilies.org', 'www.efloras.org', 'wcsp.science.kew.org', 'www.rhs.org', 'www.borealforest.org', 'biodiversitylibrary.org', 'www.rhs.org', 'wcsp.science.kew.org', 'www.esa.org', 'www.rhs.org', 'www.rhs.org', 'www.aspcapro.org', 'www.rhs.org', 'www.rhs.org', 'www.rhs.org', 'www.rhs.org', 'www.rhs.org', ['育種学雑誌 breeding science '], ['molecular phylogenetics and evolution'], ['plant systematics and evolution'], ['frontiers in plant science '], ['plant science '], ['j. am. vet. med. assoc. '], ['theoretical and applied genetics '], ['育種学雑誌 breeding science '], ['topics in companion animal medicine'], ['plant systematics and evolution ']]",73421,Allow all users (no expiry set),86619,19 August 2002,Karen Johnson ,1868,0,2002-08-19,2002-08,2002
293,293,Tamils,https://en.wikipedia.org/wiki/Tamils,187,11,"['10.2307/3516775', '10.2307/2053272', '10.2307/3516448', '10.1080/09557570701828592', '10.2307/2659023', '10.1080/01436590600850434', '10.1525/ae.1975.2.1.02a00100', '10.1353/fta.0.0031', '10.2307/2053325', '10.1086/462931', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None]","[['social scientist '], [' the journal of asian studies '], ['social scientist '], ['[[cambridge review of international affairs'], ['the journal of asian studies '], ['[[third world quarterly'], ['american ethnologist '], ['  future anterior '], ['the journal of asian studies'], ['history of religions']]",9,8,0,32,0,1,126,0.0481283422459893,0.0427807486631016,0.1711229946524064,0.058823529411764705,0.0,0.1497326203208556,10,"['www.statistics.gov', 'www.statistics.gov', 'censusindia.gov', 'censusindia.gov', 'www.singstat.gov', 'www.singstat.gov', 'censusindia.gov', 'statistics.gov', 'www.flonnet.com', 'books.google.com', 'www.britannica.com', 'www.britannica.com', 'www.hindu.com', 'www.hindustantimes.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.flonnet.com', 'books.google.com', 'newstodaynet.com', 'books.google.com', 'tamilnadu.com', 'www.hindu.com', 'www.business-standard.com', 'www.bnaiyer.com', 'www.thehindu.com', 'eelavar.com', 'gateway.proquest.com', 'www.hindu.com', 'books.google.com', 'travel.nytimes.com', 'www.flonnet.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.intamm.com', 'www.hindu.com', 'www.thenews.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'www.hrw.org', 'www.royalacademy.org', 'www.uthr.org', 'heritagetoronto.org', 'statsmauritius.govmu.org', 'www.tamilvu.org', 'tamilnation.org', 'murugan.org', 'sports.indiapress.org', ['social scientist '], [' the journal of asian studies '], ['social scientist '], ['[[cambridge review of international affairs'], ['the journal of asian studies '], ['[[third world quarterly'], ['american ethnologist '], ['  future anterior '], ['the journal of asian studies'], ['history of religions']]",300548,Allow all users (no expiry set),108811,20 August 2003,Graculus ,6225,28,2003-08-20,2003-08,2003
294,294,South India,https://en.wikipedia.org/wiki/South_India,320,9,"['10.1525/as.2002.42.5.733', '10.1080/14672715.1991.10413152', '10.1023/b:popu.0000020882.29684.8e', None, '10.1177/006996677601000202', '10.2307/3520429', '10.1038/35002501', None, None, None, '19001685', None, None, '10706275', None, None, None, None, None, None, None]","[['[[asian survey', '[[university of california press'], ['bulletin of concerned asian scholars', 'committee of concerned asian scholars'], ['population research and policy review'], ['the indian journal of medical research', 'council of social development'], ['contributions to indian sociology'], ['social scientist'], ['nature']]",16,52,0,104,0,0,139,0.05,0.1625,0.325,0.028125,0.0,0.240625,7,"['www.indianrail.gov', 'www.cia.gov', 'www.censusindia.gov', 'www.telangana.gov', 'www.telangana.gov', 'www.scr.indianrailways.gov', 'india.gov', 'www.censusindia.gov', 'censusindia.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'www.wii.gov', 'www.telangana.gov', 'www.ap.gov', 'tourism.gov', 'www.indiabudget.gov', 'www.indianrailways.gov', 'www.tnsericulture.gov', 'lcweb2.loc.gov', 'business.gov', 'www.indianrailways.gov', 'www.sr.indianrailways.gov', 'censusindia.gov', 'apsrtc.gov', 'iced.cag.gov', 'www.indianrailways.gov', 'data.gov', 'mohua.gov', 'www.tn.gov', 'www.censusindia.gov', 'knowindia.gov', 'www.sr.indianrailways.gov', 'www.kerala.gov', 'www.karnataka.gov', 'www.sr.indianrailways.gov', 'www.portal.gsi.gov', 'www.sr.indianrailways.gov', 'www.scr.indianrailways.gov', 'www.ap.gov', 'idukki.gov', 'www.imd.gov', 'knowindia.gov', 'knowindia.gov', 'www.censusindia.gov', 'www.sr.indianrailways.gov', 'censusindia.gov', 'www.sr.indianrailways.gov', 'www.censusindia.gov', 'knowindia.gov', 'www.imdchennai.gov', 'oceanservice.noaa.gov', 'data.gov', 'tamilnadu.com', 'www.britannica.com', 'timesofindia.indiatimes.com', 'www.hindu.com', 'www.sanctuaryasia.com', 'books.google.com', 'www.thehindu.com', 'www.thehindu.com', 'www.gefeg.com', 'www.britannica.com', 'www.thehindu.com', 'www.britannica.com', 'www.ndtv.com', 'www.oneindia.com', 'www.thehindubusinessline.com', 'articles.economictimes.indiatimes.com', 'www.deccanchronicle.com', 'www.hindu.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.hindu.com', 'mobiletoi.timesofindia.com', 'www.britannica.com', 'books.google.com', 'tamilnadu.com', 'articles.timesofindia.indiatimes.com', 'www.thehindu.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'www.rediff.com', 'articles.timesofindia.indiatimes.com', 'www.languageinindia.com', 'books.google.com', 'www.ibtimes.com', 'www.hindu.com', 'www.iskconhighertaste.com', 'www.britannica.com', 'www.thehindu.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'www.railtourismindia.com', 'www.britannica.com', 'www.sciencedaily.com', 'www.dnaindia.com', 'books.google.com', 'www.oxforddictionaries.com', 'www.indiatimes.com', 'archives.deccanchronicle.com', 'www.thehindu.com', 'books.google.com', 'www.thenationalnews.com', 'www.thenewsminute.com', 'www.lonelyplanet.com', 'timesofindia.indiatimes.com', 'www.oneindia.com', 'outlookindia.com', 'books.google.com', 'www.business-standard.com', 'www.deccanchronicle.com', 'www.citiindia.com', 'www.britannica.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'books.google.com', 'www.nationalgeographic.com', 'www.hindu.com', 'www.hindu.com', 'www.thehindu.com', 'www.hindu.com', 'www.britannica.com', 'www.thehindu.com', 'www.telegraphindia.com', 'indianrlys.wordpress.com', 'food.ndtv.com', 'www.resourceinvestor.com', 'www.citiindia.com', 'www.hinduonnet.com', 'www.tribuneindia.com', 'archive.financialexpress.com', 'mobiletoi.timesofindia.com', 'blogs.timesofindia.indiatimes.com', 'www.worldatlas.com', 'www.languageinindia.com', 'www.outlookindia.com', 'www.thehindu.com', 'www.indianexpress.com', 'books.google.com', 'www.firstpost.com', 'www.andhrabulletin.com', 'books.google.com', 'www.thehindu.com', 'outlookindia.com', 'query.nytimes.com', 'www.deccanchronicle.com', 'edition.cnn.com', 'www.thehindu.com', 'www.britannica.com', 'www.nytimes.com', 'www.britannica.com', 'www.keralartc.com', 'www.dnaindia.com', 'www.in.undp.org', 'www.filmfed.org', 'www.gefweb.org', 'faostat.fao.org', 'whc.unesco.org', 'www.iso.org', 'www.nhai.org', 'theinternationaljournal.org', 'www.nhai.org', 'indiaenvironmentportal.org', 'www.icrier.org', 'www.filmfed.org', 'www.un.org', 'faostat.fao.org', 'cato.org', 'www.panda.org', ['[[asian survey', '[[university of california press'], ['bulletin of concerned asian scholars', 'committee of concerned asian scholars'], ['population research and policy review'], ['the indian journal of medical research', 'council of social development'], ['contributions to indian sociology'], ['social scientist'], ['nature']]",678583,Allow all users (no expiry set),164301,25 May 2004,Robin klein ,5995,28,2004-05-25,2004-05,2004
295,295,Punjabis,https://en.wikipedia.org/wiki/Punjabis,149,3,"['10.1086/346068', '10.1093/jaarel/lix.2.339', '10.1017/s0021911808001204', '12536373', None, None, '379225', None, None]","[[' am. j. hum. genet. '], ['journal of the american academy of religion'], ['journal of asian studies']]",10,18,0,48,0,0,70,0.06711409395973154,0.12080536912751678,0.3221476510067114,0.020134228187919462,0.0,0.2080536912751678,3,"['www.stats.gov', 'censusindia.gov', 'statpak.gov', 'www.cia.gov', 'censusindia.gov', '2.census.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'www.pbs.gov', 'www.abs.gov', 'www.pbs.gov', 'www.cia.gov', 'www.censusindia.gov', 'www.pbs.gov', 'www.pbs.gov', 'www.censusindia.gov', 'pwd.punjab.gov', 'www.censusindia.gov', 'www.youtube.com', 'm.indiatvnews.com', 'books.google.com', 'krysstal.com', 'www.britannica.com', 'timesofindia.indiatimes.com', 'exoticindiaart.com', 'books.google.com', 'www.vahrehvah.com', 'thesikhencyclopedia.com', 'books.google.com', 'books.google.com', 'indianexpress.com', 'global.oup.com', 'softserv-intl.com', 'books.google.com', 'books.google.com', 'books.google.com', 'orientalarchitecture.com', 'timesofindia.indiatimes.com', 'books.google.com', 'padfield.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.phoenixnewtimes.com', 'ethnologue.com', 'exoticindiaart.com', 'books.google.com', 'sgr.sagepub.com', 'books.google.com', 'books.google.com', 'books.google.com', 'harappa.com', 'ethnologue.com', 'in.reuters.com', 'tribuneindia.com', 'wildfiregames.com', 'books.google.com', 'apnorg.com', 'books.google.com', 'worldatlas.com', 'books.google.com', 'articles.latimes.com', 'www.britannica.com', 'www.encyclopedia.com', 'harappa.com', 'books.google.com', 'livius.org', 'www.sikhcoalition.org', 'alislam.org', 'oecd.org', 'hrisouthasian.org', 'www.unhcr.org', 'www.oecd.org', 'unstats.un.org', 'livius.org', 'sikhs.org', [' am. j. hum. genet. '], ['journal of the american academy of religion'], ['journal of asian studies']]",583048,Require administrator access (no expiry set),86938,7 April 2004,Harisingh ,6044,22,2004-04-07,2004-04,2004
296,296,Punjabi culture,https://en.wikipedia.org/wiki/Punjabi_culture,9,0,[],[],1,0,0,7,0,0,1,0.1111111111111111,0.0,0.7777777777777778,0.0,0.0,0.1111111111111111,0,"['encyclopedia.com', 'indianexpress.com', 'omniglot.com', 'www.tribuneindia.com', 'newseastwest.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'ich.unesco.org']",6237447,Allow all users (no expiry set),11671,3 August 2006,James smith2 ,721,0,2006-08-03,2006-08,2006
297,297,Budapest,https://en.wikipedia.org/wiki/Budapest,280,1,"['10.2307/901850', None, None]","[['studia musicologica academiae scientiarum hungaricae ', 'akadémiai kiadó']]",18,13,0,98,0,0,150,0.06428571428571428,0.04642857142857143,0.35,0.0035714285714285713,0.0,0.11428571428571428,1,"['mfa.gov', 'trove.nla.gov', 'www.nyc.gov', 'www.nyc.gov', 'www.mfa.gov', 'www.ebeijing.gov', 'www.hipo.gov', 'trove.nla.gov', 'www.mfa.gov', 'www.nyc.gov', 'www.tel-aviv.gov', 'trove.nla.gov', 'www.census.gov', 'www.nytimes.com', 'budapestbylocals.com', 'foursquare.com', 'books.google.com', 'en.com', 'www.weather-atlas.com', 'www.fia.com', 'worldpopulationreview.com', 'www.shanghairanking.com', 'backyardgardener.com', 'operabal.com', 'books.google.com', 'euromonitor.typepad.com', 'lovelybudapest.com', 'www.bbc.com', 'www.mastercard.com', 'greatistanbul.com', 'budapest.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'innovation-cities.com', 'railwaygazette.com', 'budapest-card.com', 'www.britannica.com', 'guides.travelchannel.com', 'www.euromonitor.com', 'www.economistinsights.com', 'books.google.com', 'www.cee.siemens.com', 'books.google.com', 'www.britannica.com', 'www.britannica.com', 'www.shapedscape.com', 'www.smh.com', 'books.google.com', 'www.nytimes.com', 'goworldtravel.com', 'www.mastercard.com', 'www.euromonitor.com', 'bigseventravel.com', 'books.google.com', 'buecher.hagalil.com', 'climatemps.com', 'canadianaviationnews.wordpress.com', 'www.com', 'www.hurriyet.com', 'welovebudapest.com', 'books.google.com', 'cruise-profi.com', 'budapestarchitect.com', 'dinitrandu.com', 'books.google.com', 'books.google.com', 'www.gptoday.com', 'www.frommers.com', 'foodbycountry.com', 'www.fifa.com', 'encarta.msn.com', 'blog.euromonitor.com', 'money.cnn.com', 'www.thomaswhite.com', 'www.70-billion-pixels-budapest.com', 'www.plazacenters.com', 'www.pwc.com', 'pbase.com', 'www.emta.com', 'www.budpocketguide.com', 'budapest.com', 'www.lonelyplanet.com', 'books.google.com', 'www.nytimes.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'budapest.com', 'books.google.com', 'roommatesbudapest.com', 'www.bridgesofbudapest.com', 'simonsblogpark.com', 'books.google.com', 'simpletoremember.com', 'vilnius.com', 'www.timesofisrael.com', 'dailynewshungary.com', 'dailynewshungary.com', 'city-data.com', 'budapest.com', 'www.belmond.com', 'gislounge.com', 'www.citymayors.com', 'www.time.com', 'promote-cee.com', 'stay.com', 'budapestbydistrict.com', 'www.futuretravelexperience.com', 'www.britannica.com', 'lovelybudapest.com', 'whc.unesco.org', 'www.jewishvirtuallibrary.org', 'whc.unesco.org', 'cwur.org', 'gardenology.org', 'fwsistercities.org', 'whc.unesco.org', 'www.ushmm.org', 'globaldatalab.org', 'www.refworld.org', 'judapest.org', 'www.unhcr-centraleurope.org', 'www.refworld.org', 'www.imf.org', 'commons.wikimedia.org', 'whc.unesco.org', 'wwf.panda.org', 'www.imf.org', ['studia musicologica academiae scientiarum hungaricae ', 'akadémiai kiadó']]",36787,Require administrator access (no expiry set),208704,27 January 2002,Derek Ross ,6743,8,2002-01-27,2002-01,2002
298,298,Pyrénées-Orientales,https://en.wikipedia.org/wiki/Pyr%C3%A9n%C3%A9es-Orientales,11,0,[],[],1,0,0,0,0,0,10,0.09090909090909091,0.0,0.0,0.0,0.0,0.09090909090909091,0,['commons.wikimedia.org'],23455006,Allow all users (no expiry set),18095,10 February 2002,David Parker ,458,1,2002-02-10,2002-02,2002
299,299,Turkmens,https://en.wikipedia.org/wiki/Turkmens,118,9,"['10.1017/ehs.2020.11', '10.1017/ehs.2020.4', '10.1016/j.ara.2020.100177', '10.1371/journal.pone.0076748', '10.1371/journal.pone.0041252', '10.1023/a:1015262522048', '10.1038/s41586-018-0094-2', '10.1163/22105832-00702005', '10.1163/22105018-12340089', None, None, None, '24204668', '22815981', None, '29743675', None, None, None, None, None, '3799995', '3399854', None, None, None, None]","[['evolutionary human sciences ', '[[cambridge university press'], ['evolutionary human sciences ', '[[cambridge university press'], ['archaeological research in asia ', '[[elsevier'], ['plos one'], ['plos one'], ['russian journal of genetics'], ['[[nature ', '[[nature research'], ['language dynamics and change ', '[[brill publishers'], ['inner asia ', '[[brill publishers']]",10,8,0,29,0,0,62,0.0847457627118644,0.06779661016949153,0.2457627118644068,0.07627118644067797,0.0,0.2288135593220339,9,"['www.state.gov', '2001.ukrcensus.gov', 'lcweb2.loc.gov', 'www.state.gov', 'neutrality.gov', 'neutrality.gov', 'lcweb2.loc.gov', 'www.cia.gov', 'amazon.com', 'books.google.com', 'books.google.com', 'global.oup.com', 'books.google.com', 'books.google.com', 'kungrad.com', 'www.merriam-webster.com', 'asian-recipe.com', 'www.hauntedink.com', 'www.worldatlas.com', 'archive.aramcoworld.com', 'www.newscentralasia.com', 'issuu.com', 'www.google.com', 'www.turkmenkultur.com', 'books.google.com', 'zamanturkmenistan.com', 'www.ethnologue.com', 'turkmenportal.com', 'www.pavelicpapers.com', 'www.google.com', 'www.flayrah.com', 'www.ethnologue.com', 'books.google.com', 'www.routledge.com', 'books.google.com', 'www.google.com', 'www.google.com', 'zh.wikisource.org', 'zh.wikisource.org', 'www.turkmenistanembassy.org', 'doi.org', 'www.olympic.org', 'www.rferl.org', 'www.unhcr.org', 'www.rferl.org', 'www.wilsoncenter.org', 'iranicaonline.org', ['evolutionary human sciences ', '[[cambridge university press'], ['evolutionary human sciences ', '[[cambridge university press'], ['archaeological research in asia ', '[[elsevier'], ['plos one'], ['plos one'], ['russian journal of genetics'], ['[[nature ', '[[nature research'], ['language dynamics and change ', '[[brill publishers'], ['inner asia ', '[[brill publishers']]",1100924,Allow all users (no expiry set),76600,25 October 2004,4.63.191.85 ,1913,7,2004-10-25,2004-10,2004
300,300,Mozambique,https://en.wikipedia.org/wiki/Mozambique,146,8,"['10.1353/port.2004.0001', '10.1371/journal.pone.0198941', '10.4000/poldev.78', '10.1057/palgrave.fp.8200087', '10.1038/s41467-020-19493-3', '10.12987/yale/9780300109009.003.0005', '10.1017/s0003598x00047876', '10.1016/s0277-9536(02)00068-0', None, '29902271', None, None, '33293507', None, None, '12560007', None, '6002040', None, None, '7723057', None, None, None]","[['portuguese studies '], ['plos one'], ['international development policy '], ['french politics'], ['nature communications'], ['yale university press '], ['antiquity'], ['social science ']]",23,17,0,52,0,3,43,0.15753424657534246,0.11643835616438356,0.3561643835616438,0.0547945205479452,0.0,0.3287671232876712,8,"['www.dfid.gov', 'www.cia.gov', '2009-2017.state.gov', 'www.ine.gov', 'www.state.gov', '2009-2017.state.gov', 'state.gov', 'www.ine.gov', 'cia.gov', 'www.ine.gov', 'www.state.gov', 'dgarq.gov', 'cia.gov', '2009-2017.state.gov', 'maputo.usembassy.gov', 'ine.gov', 'www.ine.gov', 'www.greatadventuresafaris.com', 'www.afrol.com', 'www.glaenergy.com', 'www.economist.com', 'allafrica.com', 'www.bookofdaystales.com', 'www.bbc.com', 'www.irishtimes.com', 'www.youtube.com', 'www.nytimes.com', 'www.railwaygazette.com', 'allafrica.com', 'www.google.com', 'www.britannica.com', 'www.nytimes.com', 'www.business-anti-corruption.com', 'mondediplo.com', 'www.aljazeera.com', 'www.nytimes.com', 'constructionreviewonline.com', 'books.google.com', 'www.glaenergy.com', 'www.britannica.com', 'www.britannica.com', 'www.bbc.com', 'theempire.com', 'www.measuredhs.com', 'www.nytimes.com', 'www.britannica.com', 'www.indiablooms.com', 'news.com', 'apnews.com', 'books.google.com', 'foreignpolicy.com', 'forward.com', 'books.google.com', 'books.google.com', 'dhsprogram.com', 'allafrica.com', 'www.thehindubusinessline.com', 'books.google.com', 'www.news24.com', 'www.bbc.com', 'www.reuters.com', 'books.google.com', 'www.news24.com', 'www.britannica.com', 'www.bbc.com', 'www.bbc.com', 'www.dw.com', 'www.time.com', 'www.nytimes.com', 'unaids.org', 'databank.worldbank.org', 'seedtracker.org', 'journals.openedition.org', 'diocesedetete.org', 'www.ibe.unesco.org', 'ifad.org', 'hdrstats.undp.org', 'www.eisa.org', 'data.uis.unesco.org', 'communistcrimes.org', 'www.imf.org', 'moumethodist.org', 'mormonnewsroom.org', 'www.globalsecurity.org', 'www.poptel.org', 'hdr.undp.org', 'www.sahistory.org', 'communistcrimes.org', 'cpj.org', 'data.worldbank.org', 'www.content.eisa.org', 'www.unfpa.org', ['portuguese studies '], ['plos one'], ['international development policy '], ['french politics'], ['nature communications'], ['yale university press '], ['antiquity'], ['social science ']]",19301,Require administrator access (no expiry set),135982,23 May 2001,KoyaanisQatsi ,4330,8,2001-05-23,2001-05,2001
301,301,Elâzığ,https://en.wikipedia.org/wiki/El%C3%A2z%C4%B1%C4%9F,34,1,"['10.31826/hug-2020-230110', None, None]",[['hugoye']],5,4,0,9,0,0,15,0.14705882352941177,0.11764705882352941,0.2647058823529412,0.029411764705882353,0.0,0.29411764705882354,1,"['www.mgm.gov', 'kultur.gov', 'kultur.gov', 'www.dhmi.gov', 'www.world-airport-codes.com', 'haberturk.com', 'firatuniversitesi.medyasoftdigital.com', 'www.google.com', 'books.google.com', 'bilgilersitesi.com', 'books.google.com', 'en.milligazete.com', 'www.turkeyforyou.com', 'www.wdl.org', 'www.wdl.org', 'www.wdl.org', 'atonet.org', 'soc-wus.org', ['hugoye']]",2341852,Allow all users (no expiry set),30036,30 July 2005,63.98.108.24 ,1076,2,2005-07-30,2005-07,2005
302,302,Culture of Slovakia,https://en.wikipedia.org/wiki/Culture_of_Slovakia,15,0,[],[],1,0,0,4,0,0,10,0.06666666666666667,0.0,0.26666666666666666,0.0,0.0,0.06666666666666667,0,"['slovakiasite.com', 'books.google.com', 'iihf.com', 'iihf.com', 'whc.unesco.org']",11661795,Allow all users (no expiry set),16275,8 June 2007,Dr. Blofeld ,92,0,2007-06-08,2007-06,2007
303,303,"Phoenix, Arizona","https://en.wikipedia.org/wiki/Phoenix,_Arizona",355,5,"['10.1017/s0898030609090058', '10.1080/00431672.2019.1659034', None, '10.1016/j.wneu.2010.07.011', '10.5194/hess-11-1633-2007', None, None, '24979972', '21299987', None, None, None, None, None, None]","[['journal of policy history '], ['[[weatherwise'], ['national vital statistics reports ', 'cdc'], ['world neurosurgery '], ['hydrology and earth system sciences']]",45,65,0,175,0,1,65,0.1267605633802817,0.18309859154929578,0.49295774647887325,0.014084507042253521,0.0,0.323943661971831,5,"['scottsdaleaz.gov', 'www.phoenix.gov', 'www.phoenix.gov', 'geonames.usgs.gov', 'www.azleg.gov', 'www.srpmic-nsn.gov', 'www.srpmic-nsn.gov', 'www.azmag.gov', 'focus.nps.gov', 'quickfacts.census.gov', 'chroniclingamerica.loc.gov', 'www.census.gov', 'factfinder.census.gov', 'www.archives.gov', 'www.maricopa.gov', 'www.census.gov', 'www.tonation-nsn.gov', 'www.azenergy.gov', 'azmemory.azlibrary.gov', 'azsos.gov', 'quickfacts.census.gov', 'www.wrh.noaa.gov', 'w2.weather.gov', 'www.bop.gov', 'www.ade.az.gov', 'www.phoenix.gov', 'apps.bea.gov', 'census.gov', 'www.azdot.gov', 'azmemory.azlibrary.gov', 'www.azgfd.gov', 'www.census.gov', 'www.phoenix.gov', 'www.ucrdatatool.gov', 'phoenix.gov', 'www.phoenix.gov', 'www.maricopa.gov', 'factfinder.census.gov', 'www.census.gov', 'www.fbi.gov', 'geonames.usgs.gov', 'www.phoenix.gov', 'nps.gov', 'factfinder.census.gov', 'www.census.gov', 'www.gsa.gov', 'factfinder.census.gov', 'www.maricopa.gov', 'phoenix.gov', 'glorecords.blm.gov', 'factfinder.census.gov', 'www.phoenix.gov', 'www.fhwa.dot.gov', 'quickfacts.census.gov', 'www.bls.gov', 'www.census.gov', 'www2.census.gov', 'tempe.gov', 'www.bls.gov', 'www.azd.uscourts.gov', 'www.census.gov', 'jphxprd.phoenix.gov', 'factfinder.census.gov', 'www.phoenix.gov', 'geonames.usgs.gov', 'mirror-pole.com', 'www.desertusa.com', 'azbigmedia.com', 'www.tucsonsentinel.com', 'metrophoenixinvestmentproperties.listinglab.com', 'books.google.com', 'books.google.com', 'www.bizjournals.com', 'nascar.com', 'www.earlychildhoodeducationzone.com', 'www.azcentral.com', 'theculturetrip.com', 'www.srpnet.com', 'phoenix-theater.com', 'www.azcentral.com', 'cronkitenewsonline.com', 'www.nba.com', 'www.nba.com', 'www.emporis.com', 'www.marketwatch.com', 'azcentral.com', 'www.skyharbor.com', 'azheart.com', 'farmersalmanac.com', 'www.888notheft.com', 'www.smartcitiesdive.com', 'www.history.com', 'health.usnews.com', 'skyharbor.com', 'newgeography.com', 'www.amtrakconnectsus.com', 'discoverphoenix.com', 'www.azcentral.com', 'emporis.com', 'jdbaseball.com', 'www.businessinsider.com', 'www.salon.com', 'www.azcentral.com', 'www.azigg.com', 'www.azcentral.com', 'www.economist.com', 'visitphoenix.com', 'usatoday30.usatoday.com', 'www.mesa-air.com', 'azcentral.com', 'worldpopulationreview.com', 'health.usnews.com', 'www.nba.com', 'www.wnba.com', 'azenergy.com', 'wateruseitwisely.com', 'www.weather-us.com', 'www.nytimes.com', 'mlb.mlb.com', 'www.azcentral.com', 'fcx.com', 'www.marketingcharts.com', 'www.azstarnet.com', 'www.historicphoenix.com', 'www.cbs5az.com', 'www.smartcitiesdive.com', 'www.emporis.com', 'www.wnba.com', 'health.usnews.com', 'wnba.com', 'www.drugaddictiontreatment.com', 'azfamily.com', 'www.wsj.com', 'azcentral.com', 'www.azcentral.com', 'www.barriozona.com', 'aerospace.honeywell.com', 'health.usnews.com', 'www.azcentral.com', 'www.archdaily.com', 'www.washingtonpost.com', 'www.usnpl.com', 'bleacherreport.com', 'www.nfl.com', 'skyscraperpage.com', 'www.cnn.com', 'www.emporis.com', 'www.phoenixchamber.com', 'www.azcentral.com', 'phoenixasap.com', 'www.nbcnews.com', 'skyharbor.com', 'www.worldatlas.com', 'www.thearda.com', 'www.azcentral.com', 'archive.azcentral.com', 'www.visitphoenix.com', 'skyharbor.com', 'wmphoenixopen.com', 'health.usnews.com', 'www.foxnews.com', 'www.eastvalleytribune.com', 'www.asugammage.com', 'www.discoverphoenixarizona.com', 'phoenix.about.com', 'www.foxnews.com', 'history.com', 'origin.nba.com', 'phoenix.about.com', 'www.arizonaedventures.com', 'frontdoorsnews.com', 'www.phoenixnewtimes.com', 'www.nba.com', 'books.google.com', 'www.azcentral.com', 'www.azcentral.com', 'history.com', 'www.azcentral.com', 'sportsecyclopedia.com', 'www.lpgafounderscup.com', 'books.google.com', 'www.mnn.com', 'www.nfl.com', 'locations.greyhound.com', 'ezinemark.com', 'www.phoenixsnakeremoval.com', 'www.forbes.com', 'books.google.com', 'www.azcentral.com', 'stockyardssteakhouse.com', 'www.arizonascots.com', 'www.historycentral.com', 'www.azcentral.com', 'www.nba.com', 'www.azcentral.com', 'about.com', 'www.residentialarchitect.com', 'www.cap-az.com', 'www.slamonline.com', 'phoenix.about.com', 'www.macayo.com', 'skyharbor.com', 'www.azcardinals.com', 'ktar.com', 'phoenix-az.knoji.com', 'phoenixraceway.com', 'health.usnews.com', 'queencreekindependent.com', 'www.azcentral.com', 'azcentral.com', 'money.cnn.com', 'abcnews.go.com', 'content.time.com', 'baseball-reference.com', 'visitphoenix.com', 'about.com', 'phoenix.about.com', 'www.huffingtonpost.com', 'azcentral.com', 'ratings.radio-online.com', 'www.nba.com', 'www.accessgenealogy.com', 'www.abc15.com', 'www.phoenixnewtimes.com', 'www.discoverphoenixarizona.com', 'coyotes.nhl.com', 'usatoday30.usatoday.com', 'nascar.com', 'texaseagle.com', 'phoenixrestaurants.com', 'www.jcl.com', 'intel.com', 'www.residentialarchitect.com', 'www.bizjournals.com', 'www.arizonaguide.com', 'www.phoenixnewtimes.com', 'www.accessgenealogy.com', 'www.history.com', 'www.baseball-almanac.com', 'www.bannerhealth.com', 'www.lung.org', 'www.transportation-finance.org', 'phxart.org', 'phoenixzoo.org', 'arizonaexperience.org', 'cloud.tpl.org', 'www.itheatreaz.org', 'trainweb.org', 'www.valleymetro.org', 'ballotpedia.org', 'www.phoenixsistercities.org', 'www.dbg.org', 'azfo.org', 'www.mcso.org', 'heard.org', 'www.lung.org', 'www.phoenixsistercities.org', 'www.diocesephoenix.org', 'desertmuseum.org', 'azchallenger.org', 'www.gilariver.org', 'www.researchhistory.org', 'www.pewresearch.org', 'www.ccrh.org', 'www.mayoclinic.org', 'www.arizonaexperience.org', 'www.pewforum.org', 'www.sanxaviermission.org', 'arizonahistoricalsociety.org', 'fiestabowl.org', 'fiestabowl.org', 'herbergertheater.org', 'trainweb.org', 'azta.org', 'estrellawar.org', 'www.nicb.org', 'phoenixopera.org', 'mirandawarning.org', 'phoenixsistercities.org', 'summitpost.org', 'jstor.org', 'www.america2050.org', 'www.desertmuseum.org', 'davesredistricting.org', 'www.mayoclinic.org', ['journal of policy history '], ['[[weatherwise'], ['national vital statistics reports ', 'cdc'], ['world neurosurgery '], ['hydrology and earth system sciences']]",49121,Allow all users (no expiry set),210227,15 April 2002,Jeronimo ,7977,25,2002-04-15,2002-04,2002
304,304,Mykonos,https://en.wikipedia.org/wiki/Mykonos,40,1,"['10.1080/19443994.2012.714603', None, None]",[['desalination and water treatment']],0,0,0,26,0,0,13,0.0,0.0,0.65,0.025,0.0,0.025,1,"['www.inmykonos.com', 'books.google.com', 'www.inmykonos.com', 'www.collinsdictionary.com', 'www.inmykonos.com', 'www.inmykonos.com', 'www.inmykonos.com', 'www.inmykonos.com', 'article.wn.com', 'www.inmykonos.com', 'www.inmykonos.com', 'books.google.com', 'travelwideworld.com', 'www.inmykonos.com', 'www.inmykonos.com', 'www.inmykonos.com', 'www.inmykonos.com', 'www.mykonos-web.com', 'greeka.com', 'www.inmykonos.com', 'www.inmykonos.com', 'www.mykonos-airport.com', 'www.inmykonos.com', 'www.inmykonos.com', 'www.inmykonos.com', 'www.mykonos-accommodation.com', ['desalination and water treatment']]",490946,Allow all users (no expiry set),31679,27 February 2004,Adam Bishop ,1710,3,2004-02-27,2004-02,2004
305,305,Buryats,https://en.wikipedia.org/wiki/Buryats,48,18,"['10.1002/ajhb.23194', '10.1163/000000009793066596', '10.1134/s1022795413110082', 'abs/10.1080/10758216.2015.1057040', '10.1007/s100380050015', '10.1163/146481700793647931', '10.1007/s10038-005-0322-0', '10.1111/j.1469-1809.2010.00601.x', '10.1086/soutjanth.10.3.3629134', '10.1046/j.1529-8817.2003.00127.x', '10.1007/s00439-005-0076-y', None, '10.2307/2696979', '10.1186/2041-2223-2-10', '10.1086/522933', '10.1038/s41586-021-03336-2', '10.1086/710574', '10.1086/338457', '30408262', None, None, None, '10721667', None, '16328082', '20726964', None, '15638829', '16261343', '11236866', None, '21463511', '17924343', None, None, '11731934', None, None, None, None, None, None, None, None, None, '3905771', None, None, None, '3087676', '2265662', None, None, '384887']","[['american journal of human biology '], ['inner asia '], ['russian journal of genetics '], ['problems of post-communism '], ['journal of human genetics '], ['inner asia '], ['journal of human genetics '], ['annals of human genetics '], ['southwestern journal of anthropology '], ['annals of human genetics '], ['human genetics '], ['human biology '], ['slavic review '], ['investigative genetics '], ['the american journal of human genetics '], ['nature'], ['[[history of religions ', '[[university of chicago press'], ['the american journal of human genetics ']]",4,0,0,4,0,0,22,0.08333333333333333,0.0,0.08333333333333333,0.375,0.0,0.4583333333333333,18,"['ethnologue.com', 'jsbednet.com', 'brill.com', 'www.yfull.com', 'www.culturalsurvival.org', 'www.unspecial.org', 'sreda.org', 'www.unesco.org', ['american journal of human biology '], ['inner asia '], ['russian journal of genetics '], ['problems of post-communism '], ['journal of human genetics '], ['inner asia '], ['journal of human genetics '], ['annals of human genetics '], ['southwestern journal of anthropology '], ['annals of human genetics '], ['human genetics '], ['human biology '], ['slavic review '], ['investigative genetics '], ['the american journal of human genetics '], ['nature'], ['[[history of religions ', '[[university of chicago press'], ['the american journal of human genetics ']]",57701,Allow all users (no expiry set),48881,17 June 2002,Peterlin~enwiki ,664,8,2002-06-17,2002-06,2002
306,306,Culture of Japan,https://en.wikipedia.org/wiki/Culture_of_Japan,63,5,"['10.1126/sciadv.abh2419', '10.2307/3773912', '10.2307/3112093', '10.1038/jhg.2016.110', '10.1093/jdh/8.3.215', '34533991', None, None, '27581845', None, '8448447', None, None, '5285490', None]","[['science advances '], [' ethnology'], [' the business history review'], [' journal of human genetics'], [' journal of design history']]",8,0,0,18,0,1,31,0.12698412698412698,0.0,0.2857142857142857,0.07936507936507936,0.0,0.20634920634920634,5,"['public.oed.com', 'public.oed.com', 'www.asahi.com', 'books.google.com', 'www.omniglot.com', 'nippon.com', 'www.asianweek.com', 'japan-and-mexico-meet.tumblr.com', 'urushi-joboji.com', 'theconversation.com', 'www.usnews.com', 'livescience.com', 'www.reuters.com', 'www.tokyohive.com', 'qz.com', 'blog.ratestogo.com', 'www.channelnewsasia.com', 'www.forbes.com', 'libmma.contentdm.oclc.org', 'japanfocus.org', 'dcaj.org', 'web-japan.org', 'web-japan.org', 'web-japan.org', 'www.sljfaq.org', 'www.sljfaq.org', ['science advances '], [' ethnology'], [' the business history review'], [' journal of human genetics'], [' journal of design history']]",167104,Allow all users (no expiry set),56633,9 January 2003,TakuyaMurata ,4870,13,2003-01-09,2003-01,2003
307,307,Basques,https://en.wikipedia.org/wiki/Basques,72,20,"['10.1073/pnas.1509851112', '10.1186/1471-2164-7-124', '10.1016/j.ajhg.2012.01.002', '10.1371/journal.pbio.1000285', '10.1126/science.290.5494.1155', '10.1038/s41598-021-84915-1', '10.1126/science.aav4040', '10.1038/ejhg.2010.146', '10.1038/sj.ejhg.5201482', '10.1038/s41598-017-07710-x', '10.1038/s41467-018-08272-w', '10.1017/s0020859005002087', '10.1093/molbev/msi185', '10.1126/science.1153717', '10.1016/j.ympev.2006.11.030', '10.1007/s00439-010-0833-4', '10.1371/journal.pone.0021592', '10.1093/molbev/msh135', '10.1126/science.aax3372', '10.1080/713683438', '26351665', '16719915', '22365151', '20087410', '11073453', '33692401', '30872528', '20736979', '16094307', '28779148', '30710075', None, '15944443', '18292342', '17275346', '20443121', '21720564', '15044595', None, None, '4586848', '1523212', '3309182', '2799514', None, '7970938', '6436108', '3039512', None, '5544771', '6358624', None, None, None, None, None, '3123369', None, None, None]","[['proceedings of the national academy of sciences'], ['bmc genomics'], ['the american journal of human genetics'], [' [[plos biology', ' [[public library of science'], ['sciencemag.org ', 'science '], ['scientific reports'], ['science'], ['european journal of human genetics', 'springer nature'], ['european journal of human genetics ', 'springer nature '], ['[[scientific reports'], ['nature communications'], ['international review of social history'], ['molecular biology and evolution', 'oxford university press'], ['science'], ['mol. phylogenet. evol. '], ['human genetics'], ['plos one', 'public library of science'], ['molecular biology and evolution', 'oxford university press'], ['[[science '], ['journal of spanish cultural studies ']]",7,1,0,13,0,0,31,0.09722222222222222,0.013888888888888888,0.18055555555555555,0.2777777777777778,0.0,0.3888888888888889,20,"['www.census.gov', 'books.google.com', 'kids.britannica.com', 'books.google.com', 'www.nationalgeographic.com', 'www.oxfordreference.com', 'maire-info.com', 'www.bbc.com', 'www.noticiasdenavarra.com', 'eitb24.com', 'books.google.com', 'www.eitb.com', 'books.google.com', 'the-scientist.com', 'euskomedia.org', 'www.americamagazine.org', 'basqueed.org', 'phys.org', '5d_anthropological_genetics_th(bookzz.org', '5d_anthropological_genetics_th(bookzz.org', 'filosofia.org', ['proceedings of the national academy of sciences'], ['bmc genomics'], ['the american journal of human genetics'], [' [[plos biology', ' [[public library of science'], ['sciencemag.org ', 'science '], ['scientific reports'], ['science'], ['european journal of human genetics', 'springer nature'], ['european journal of human genetics ', 'springer nature '], ['[[scientific reports'], ['nature communications'], ['international review of social history'], ['molecular biology and evolution', 'oxford university press'], ['science'], ['mol. phylogenet. evol. '], ['human genetics'], ['plos one', 'public library of science'], ['molecular biology and evolution', 'oxford university press'], ['[[science '], ['journal of spanish cultural studies ']]",4660,Allow all users (no expiry set),89465,23 November 2001,62.174.12.xxx ,3854,10,2001-11-23,2001-11,2001
308,308,Somalia,https://en.wikipedia.org/wiki/Somalia,351,18,"['10.1080/17531050903273719', '10.1016/j.quaint.2014.04.038', '10.1002/jid.1482', '10.1126/science.1078208', '10.1080/09692290701869688', '10.1007/s10437-008-9032-2', '10.1017/s0020743800063145', '10.1080/00438243.1988.9980055', '10.1525/ae.1975.2.4.02a00030', '10.1162/isec.2007.31.3.74', '10.1186/1476-072x-9-45', None, '10.1007/bf01540131', '10.2307/217389', '10.1093/biosci/bix014', '10.2307/2840281', '10.3406/ethio.1976.1157', '10.1111/j.1740-9713.2014.00717.x', None, None, None, '12714734', None, None, None, '16470993', None, None, '20840751', '17903054', None, None, '28608869', None, None, None, None, None, None, None, None, None, None, None, None, None, '2949749', None, None, None, '5451287', None, None, None]","[['journal of eastern african studies'], ['quaternary international'], ['journal of international development'], [' science '], ['review of international political economy'], ['african archaeological review'], ['international journal of middle east studies'], ['world archaeology'], ['american ethnologist '], ['international security'], ['international journal of health geographics'], ['archives of iranian medicine'], [' computers and translation '], ['[[the international journal of african historical studies'], ['bioscience'], ['[[man '], ['annales d'], ['significance']]",48,11,0,113,0,2,159,0.13675213675213677,0.03133903133903134,0.32193732193732194,0.05128205128205128,0.0,0.21937321937321938,18,"['permanent.access.gpo.gov', 'lcweb2.loc.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'travel.state.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'lcweb2.loc.gov', 'education.puntlandgovt.com', 'books.google.com', 'education.puntlandgovt.com', 'www.thejakartapost.com', 'www.voanews.com', 'books.google.com', 'garoweonline.com', 'education.puntlandgovt.com', 'somaliweyn.com', 'books.google.com', 'books.google.com', 'togdheernews.com', 'www.nytimes.com', 'education.puntlandgovt.com', 'books.google.com', 'www.independent.com', 'news.xinhuanet.com', 'blogs.nationalgeographic.com', 'www.innercitypress.com', 'www.bbc.com', 'books.google.com', 'news.google.com', 'www.aljazeera.com', 'books.google.com', 'books.google.com', 'books.google.com', 'twitter.com', 'www.ethnologue.com', 'sabahionline.com', 'www.africanexecutive.com', 'www.washingtonexaminer.com', 'books.google.com', 'education.puntlandgovt.com', 'education.puntlandgovt.com', 'www.somalilandlaw.com', 'books.google.com', 'www.youtube.com', 'bartleby.com', 'books.google.com', 'garoweonline.com', 'books.google.com', 'ameinfo.com', 'www.businessweek.com', 'www.banadir.com', 'www.google.com', 'www.reuters.com', 'www.garoweonline.com', 'archive.wikiwix.com', 'www.afrol.com', 'books.google.com', 'books.google.com', 'www.flightglobal.com', 'books.google.com', 'gulfnews.com', 'books.google.com', '(ft.com', 'www.aa.com', 'www.nytimes.com', 'www.busiweek.com', 'www.bbc.com', 'www.marketwatch.com', 'www.qurbejoog.com', 'www.google.com', 'news.xinhuanet.com', 'books.google.com', 'www.nytimes.com', 'goobjoog.com', 'books.google.com', 'strategypage.com', 'dictionary.com', 'books.google.com', 'www.google.com', 'somalilandgov.com', 'www.google.com', 'www.raxanreeb.com', 'www.google.com', 'books.google.com', 'books.google.com', 'education.puntlandgovt.com', 'www.nytimes.com', 'www.somaliweyn.com', 'www.google.com', 'sabahionline.com', 'gantdaily.com', 'books.google.com', 'books.google.com', 'books.google.com', 'dastuurkeenna.com', 'www.tashiwanaag.com', 'www.britannica.com', 'www.peterleeson.com', 'buluugleey.com', 'goobjoog.com', 'education.puntlandgovt.com', 'www.somenergy.com', 'www.wsj.com', 'lexico.com', 'www.arabnews.com', 'books.google.com', 'scribd.com', 'allafrica.com', 'books.google.com', 'education.puntlandgovt.com', 'books.google.com', 'www.newyorker.com', 'books.google.com', 'blogs.ft.com', 'www.howwemadeitinafrica.com', 'sabahionline.com', 'health.puntlandgovt.com', 'www.fiba.com', 'www.waltainfo.com', 'sabahionline.com', 'unctad.org', 'data.un.org', 'www.oic-oci.org', 'globalpolicy.org', 'lettre-ulysses-award.org', 'www.diaspora-centre.org', 'somalbanca.org', 'www.crisisgroup.org', 'www.unaids.org', 'www.ri.org', 'somalia.unfpa.org', 'www.crisisgroup.org', 'www.iaea.org', 'www.care-international.org', 'www.unhcr.org', 'www.care-international.org', 'unep.org', 'www.un.org', 'unis.unvienna.org', 'www.goldmanprize.org', 'cal.org', 'meeting.physanth.org', 'www.cfr.org', 'www.lasportal.org', 'imf.org', 'somalia.unfpa.org', 'www.unhcr.org', 'www.nti.org', 'somalbanca.org', 'www.cfr.org', 'www.oic-oci.org', 'www.pewforum.org', 'amisom-au.org', 'cal.org', 'www.unfpa.org', 'afjn.org', 'www.un.org', 'www.kenyahighcomtz.org', 'data.worldbank.org', 'unpos.unmissions.org', 'www.opec.org', 'population.un.org', 'somalbanca.org', 'mepc.org', 'www.hornrelief.org', 'wes.org', 'www.reptile-database.org', 'www.elmt-relpa.org', ['journal of eastern african studies'], ['quaternary international'], ['journal of international development'], [' science '], ['review of international political economy'], ['african archaeological review'], ['international journal of middle east studies'], ['world archaeology'], ['american ethnologist '], ['international security'], ['international journal of health geographics'], ['archives of iranian medicine'], [' computers and translation '], ['[[the international journal of african historical studies'], ['bioscience'], ['[[man '], ['annales d'], ['significance']]",27358,Require administrator access (no expiry set),215073,27 May 2001,KoyaanisQatsi ,13634,27,2001-05-27,2001-05,2001
309,309,Occitania,https://en.wikipedia.org/wiki/Occitania,124,1,[],[],7,0,0,22,0,0,94,0.056451612903225805,0.0,0.1774193548387097,0.008064516129032258,0.0,0.06451612903225806,0,"['fr.dir.groups.yahoo.com', 'www.hcplive.com', 'books.google.com', 'www.paugolfclub.com', 'www.jornalet.com', 'books.google.com', 'myriamchabrun.chez.com', 'www.jornalet.com', 'www.ben-vautier.com', 'media.wix.com', 'opinion.jornalet.com', 'www.festival-douarnenez.com', 'books.google.com', 'www.lexilogos.com', 'books.google.com', 'resultados.elpais.com', 'books.google.com', 'www.elsevier.com', 'www.xarnege.com', 'books.google.com', 'books.google.com', 'www.gasconha.com', 'upload.wikimedia.org', 'upload.wikimedia.org', 'www.arkheia-revue.org', 'www.p-n-o.org', 'upload.wikimedia.org', 'www.minorityrights.org', 'www.museeprotestant.org']",1149357,Allow all users (no expiry set),108884,9 November 2004,62.147.90.102 ,1346,4,2004-11-09,2004-11,2004
310,310,Yakuts,https://en.wikipedia.org/wiki/Yakuts,60,9,"[None, '10.1017/s0041977x00005498', '10.1186/1471-2148-13-127', '10.20874/2071-0437-2018-41-2-119-127', '10.17223/15617793/407/23', '10.1371/journal.pone.0083570', '10.17516/1997-1370-2016-9-8-1822-1840', '10.1016/j.aeae.2011.08.012', '10.22162/2619-0990-2020-50-4-941-950', '18610830', None, '23782551', None, None, '24349531', None, None, None, None, None, '3695835', None, None, '3861515', None, None, None]","[['molekuliarnaia biologiia'], ['bulletin of the school of oriental and african studies'], ['bmc evolutionary biology'], ['vestnik arheologii', 'institute for humanities research and indigenous studies of the north'], ['vestnik tomskogo gosudarstvennogo universiteta', 'institute of the humanities and the indigenous peoples'], ['plos one'], ['journal of siberian federal university humanities and social sciences'], ['archaeology'], ['oriental studies', 'east siberian state institute of culture']]",1,3,0,6,0,0,41,0.016666666666666666,0.05,0.1,0.15,0.0,0.21666666666666667,9,"['data.gov', 'www.pmlp.gov', 'www.ukrcensus.gov', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.insidethenewrussia.com', 'aklyosov.home.com', 'unesdoc.unesco.org', ['molekuliarnaia biologiia'], ['bulletin of the school of oriental and african studies'], ['bmc evolutionary biology'], ['vestnik arheologii', 'institute for humanities research and indigenous studies of the north'], ['vestnik tomskogo gosudarstvennogo universiteta', 'institute of the humanities and the indigenous peoples'], ['plos one'], ['journal of siberian federal university humanities and social sciences'], ['archaeology'], ['oriental studies', 'east siberian state institute of culture']]",483558,Allow all users (no expiry set),44191,23 February 2004,Joy ,974,1,2004-02-23,2004-02,2004
311,311,Egypt,https://en.wikipedia.org/wiki/Egypt,302,3,"['10.1080/1369183x.2015.1049940', '10.1177/001654928002600202', '10.1080/13530194.2015.1102708', None, None, None, None, None, None]","[['journal of ethnic and migration studies'], ['gazette '], ['british journal of middle eastern studies']]",58,25,0,110,0,5,102,0.19205298013245034,0.08278145695364239,0.36423841059602646,0.009933774834437087,0.0,0.2847682119205298,3,"['www.capmas.gov', 'www.cia.gov', 'www.sis.gov', 'www.cia.gov', 'uscirf.gov', 'www.sis.gov', 'purl.fdlp.gov', 'capmas.gov', 'capmas.gov', 'www.egypt.gov', 'www.sis.gov', 'www.eia.gov', 'capmas.gov', 'sis.gov', 'www.sis.gov', 'webarchive.nationalarchives.gov', 'capmas.gov', '2001-2009.state.gov', '2009-2017.state.gov', 'www.america.gov', 'www.capmas.gov', 'cia.gov', 'www.sis.gov', '2009-2017.state.gov', 'capmas.gov', 'tbsjournal.com', 'www.egyptindependent.com', 'www.washingtonpost.com', 'www.dailynewsegypt.com', 'www.nytimes.com', 'www.businesstodayegypt.com', 'www.washingtonpost.com', 'www.reuters.com', 'www.dailynewsegypt.com', 'www.wsj.com', 'af.reuters.com', 'www.google.com', 'www.al-monitor.com', 'www.nytimes.com', 'www.foreignpolicy.com', 'www.wsj.com', 'www.nature.com', 'weeklystandard.com', 'gulfnews.com', 'www.dailynewsegypt.com', 'www.bbc.com', 'foreignpolicy.com', 'www.nytimes.com', 'edition.cnn.com', 'books.google.com', 'www.jpost.com', 'spaceflightnow.com', 'edition.cnn.com', 'thediplomat.com', 'books.google.com', 'www.businesstodayegypt.com', 'books.google.com', 'www.theglobeandmail.com', 'www.foreignpolicy.com', 'www.bbc.com', 'www.sfgate.com', 'weatherbase.com', 'www.bbc.com', 'www.nytimes.com', 'books.google.com', 'www.fivb.com', 'af.reuters.com', 'archive.fiba.com', 'www.ewtn.com', 'www.dw.com', 'www.nytimes.com', 'books.google.com', 'www.sciencedaily.com', 'www.nytimes.com', 'www.nytimes.com', 'www.huffingtonpost.com', 'globalsurance.com', 'books.google.com', 'indexmundi.com', 'books.google.com', 'www.chinadaily.com', 'www.aljazeera.com', 'www.youregypt.com', 'www.latimes.com', 'economist.com', 'www.dailystaregypt.com', 'thediplomat.com', 'books.google.com', 'www.washingtonpost.com', 'www.nytimes.com', 'edition.cnn.com', 'www.reuters.com', 'www.washingtonpost.com', 'melitensiawth.com', 'www.aljazeera.com', 'news.sky.com', 'books.google.com', 'www.aljazeera.com', 'www.washingtonpost.com', 'abcnews.go.com', 'www.huffingtonpost.com', 'www.nytimes.com', 'books.google.com', 'news.yahoo.com', 'www.voanews.com', 'www.bbc.com', 'books.google.com', 'www.jpost.com', 'archive.fiba.com', 'egyptianstreets.com', 'www.reuters.com', 'books.google.com', 'www.csmonitor.com', 'www.reuters.com', 'egypttoday.com', 'www.foxnews.com', 'africa.reuters.com', 'encarta.msn.com', 'books.google.com', 'www.galaxie.com', 'www.bbc.com', 'www.nytimes.com', 'www.foreignaffairs.com', 'www.egyptindependent.com', 'books.google.com', 'ameinfo.com', 'www.washingtonpost.com', 'books.google.com', 'books.google.com', 'qz.com', 'books.google.com', 'news.sky.com', 'egy-map.com', 'news.yahoo.com', 'www.aljazeera.com', 'nchregypt.org', 'foodfirst.org', 'hrw.org', 'npr.org', 'www.sesrtcic.org', 'poll2017.trust.org', 'irinnews.org', 'pewforum.org', 'hrw.org', 'imf.org', 'www.chathamhouse.org', 'irinnews.org', 'english.ahram.org', 'research.policyarchive.org', 'data.worldbank.org', 'www.worldaffairsjournal.org', 'www.jhsonline.org', 'www.pewforum.org', 'www.oecd-ilibrary.org', 'english.ahram.org', 'ancientsudan.org', 'www.worldtimelines.org', 'english.ahram.org', 'weekly.ahram.org', 'globalsecurity.org', 'www.ilo.org', 'english.ahram.org', 'www.fungal-conservation.org', 'hosted.ap.org', 'www.sesrtcic.org', 'english.ahram.org', 'www.undp-pogar.org', 'www.pewglobal.org', 'www.persecutionofahmadis.org', 'hdr.undp.org', 'pewforum.org', 'undp.org', 'www.eohr.org', 'www.pewforum.org', 'english.ahram.org', 'english.ahram.org', 'freedomhouse.org', 'fas.org', 'en.eohr.org', 'english.ahram.org', 'jcpa.org', 'www.pewglobal.org', 'english.ahram.org', 'www.freedomhouse.org', 'fidh.org', 'english.ahram.org', 'modernegypt.bibalex.org', 'marketplace.publicradio.org', 'amnesty.org', 'www.unicef.org', 'carnegie-mec.org', 'www.imf.org', 'www.pewforum.org', ['journal of ethnic and migration studies'], ['gazette '], ['british journal of middle eastern studies']]",8087628,Require administrator access (no expiry set),236708,31 October 2001,Corvus13 ,11018,20,2001-10-31,2001-10,2001
312,312,Guimarães,https://en.wikipedia.org/wiki/Guimar%C3%A3es,9,0,[],[],0,0,0,4,0,0,5,0.0,0.0,0.4444444444444444,0.0,0.0,0.0,0,"['www.imdb.com', 'portugalromano.com', 'www.nytimes.com', 'www.imdb.com']",24740448,Allow all users (no expiry set),34171,18 October 2009,TrueColour ,401,0,2009-10-18,2009-10,2009
313,313,Kuwait,https://en.wikipedia.org/wiki/Kuwait,592,21,"['10.1186/s12913-018-2960-x', '10.5334/ai.0613', '10.3109/10401239309148971', '10.1017/qua.2022.3', '10.25159/1947-9417/3435', '10.1111/aae.12145', '10.1080/13530190500281424', '10.2148/benv.40.1.101', '10.1080/13530194.2015.1102708', 'abs/10.1177/2347798920940081', '10.1111/aae.12195', '10.1002/dys.361', '10.3390/resources7030058', '10.1215/1089201x-3139815', '10.1016/s0011-9164(01)00259-4', '10.1080/00263206.2011.565143', '10.1111/aae.12190', '10.1080/14634988.2012.663706', '10.20991/allazimuth.960945', '10.1111/j.1600-0471.2007.00283.x', '29510705', None, '8348201', None, None, None, None, None, None, None, None, '18433005', None, None, None, None, None, None, None, None, '5840785', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None]","[['[[bmc health services research'], ['archaeology international'], ['annals of clinical psychiatry'], ['quaternary research'], ['education as change'], ['arabian archaeology and epigraphy'], ['british journal of middle eastern studies'], ['built environment '], ['british journal of middle eastern studies'], ['contemporary review of the middle east'], [' arabian archaeology and epigraphy'], ['dyslexia'], ['resources'], ['[[comparative studies of south asia'], ['desalination'], ['middle eastern studies'], ['arabian archaeology and epigraphy'], ['aquatic ecosystem health '], ['all azimuth'], ['jacques connan']]",108,20,0,241,0,2,200,0.18243243243243243,0.033783783783783786,0.40709459459459457,0.03547297297297297,0.0,0.2516891891891892,20,"['www.uspto.gov', 'www.cia.gov', 'aad.archives.gov', 'stat.paci.gov', 'www.cia.gov', 'earthobservatory.nasa.gov', '2009-2017.state.gov', 'stat.paci.gov', '2009-2017.state.gov', 'www.cia.gov', 'www.nasa.gov', 'www.cia.gov', 'www.csb.gov', 'earthshots.usgs.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'kdipa.gov', 'www.loc.gov', 'www.loc.gov', 'www.realwire.com', 'www.nytimes.com', 'www.bbc.com', 'books.google.com', 'hyperallergic.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.youtube.com', 'www.kuwaitbuildingshow.com', 'www.hydrocarbonprocessing.com', 'www.orbital-space.com', 'newkuwaitsummit.com', 'www.britains-smallwars.com', 'www.youtube.com', 'www.steelorbis.com', 'www.al-monitor.com', 'www.arabianbusiness.com', 'books.google.com', 'www.p2bk.com', 'arabspacenews.com', 'www.gdnonline.com', 'www.google.com', 'books.google.com', 'www.cbastudios.com', 'gulfnews.com', 'books.google.com', 'www.youtube.com', 'thearabweekly.com', 'www.iihf.com', 'books.google.com', 'books.google.com', 'www.yourmiddleeast.com', 'www.aljazeera.com', 'books.google.com', 'investvine.com', 'jacc-kw.com', 'books.google.com', 'foodsecurityindex.eiu.com', 'www.ft.com', 'www.constructionweekonline.com', 'www.thedailybeast.com', 'technology.ihs.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'arabianbusiness.com', 'www.thebusinessyear.com', 'www.thewire.com', 'gbtimes.com', 'www.theworldfolio.com', 'gulfnews.com', 'encarta.msn.com', 'search.proquest.com', 'www.bbc.com', 'cosmopolitantdaily.com', 'books.google.com', 'www.arabhealthonline.com', 'books.google.com', 'books.google.com', 'www.merriam-webster.com', 'www.arabtimesonline.com', 'books.google.com', 'www.madamasr.com', 'books.google.com', 'books.google.com', 'www.hasanews.com', 'books.google.com', 'www.birdguides.com', 'eng.alostouramagazine.com', 'www.gfmag.com', 'books.google.com', 'myartguides.com', 'books.google.com', 'al-seyassah.com', 'books.google.com', 'us.practicallaw.com', 'www.analysysmason.com', 'www.emirates247.com', 'www.worldstopexports.com', 'books.google.com', 'books.google.com', 'www.bq-magazine.com', 'thearabweekly.com', 'ameinfo.com', 'books.google.com', 'www.youtube.com', 'books.google.com', 'www.bbc.com', 'books.google.com', 'www.aljazeera.com', 'gradworks.umi.com', 'gulfnews.com', 'books.google.com', 'www.haaretz.com', 'www.zawya.com', 'www.reuters.com', 'www.ancientportsantiques.com', 'books.google.com', 'www.argusmedia.com', 'books.google.com', 'www.washingtonpost.com', 'www.epicos.com', 'www.britannica.com', 'gradworks.umi.com', 'www.xinhuanet.com', 'www.orientplanet.com', 'gradworks.umi.com', 'www.nytimes.com', 'www.khalifaqattan.com', 'advisor.museumsandheritage.com', 'www.statista.com', 'berlinarchaeology.files.wordpress.com', 'reconnectingarts.com', 'chronicle.fanack.com', 'y-oman.com', 'www.reuters.com', 'qz.com', 'www.endurosat.com', 'books.google.com', 'www.pressreader.com', 'articles.latimes.com', 'www.investopedia.com', 'www.zawya.com', 'www.arabianbusiness.com', 'www.euromoney.com', 'www.pwc.com', 'gbtimes.com', 'gulfconstructiononline.com', 'www.albawaba.com', 'books.google.com', 'books.google.com', 'www.wsj.com', 'www.google.com', 'books.google.com', 'ateliervoyage.com', 'www.orbital-space.com', 'www.tamdeen.com', 'www.hydrocarbons-technology.com', 'capkuwait.com', 'www.zawya.com', 'books.google.com', 'anba.com', 'books.google.com', 'www.icis.com', 'www.al-monitor.com', 'finance.yahoo.com', 'books.google.com', 'gulfnews.com', 'books.google.com', 'www.bloomberg.com', 'www.jadaliyya.com', 'www.al-monitor.com', 'www.oxfordbusinessgroup.com', 'www.brill.com', 'www.broadcastprome.com', 'maps.wunderground.com', 'books.google.com', 'books.google.com', 'en.oxforddictionaries.com', 'www.albawaba.com', 'books.google.com', 'alshaheedparkmuseums.com', 'research.hktdc.com', 'books.google.com', 'www.iihf.com', 'chronicle.fanack.com', 'www.bookdepository.com', 'books.google.com', 'books.google.com', 'al-seyassah.com', 'www.youtube.com', 'books.google.com', 'www.fitchratings.com', 'oxfordbusinessgroup.com', 'gulfnews.com', 'santandertrade.com', 'books.google.com', 'www.oxfordbusinessgroup.com', 'gradworks.umi.com', 'www.britannica.com', 'www.washingtonpost.com', 'articles.latimes.com', 'zinco-greenroof.com', 'www.albawaba.com', 'kipic.com', 'www.meedprojects.com', 'www.counterextremism.com', 'www.arabianbusiness.com', 'search.proquest.com', 'www.entrepreneur.com', 'www.business-anti-corruption.com', 'books.google.com', 'reconnectingarts.com', 'books.google.com', 'www.argusmedia.com', 'books.google.com', 'www.arabosounds.com', 'www.economist.com', 'www.worldpoliticsreview.com', 'www.bloomberg.com', 'books.google.com', 'www.bloomberg.com', 'books.google.com', 'arabianbusiness.com', 'books.google.com', 'www.reuters.com', 'www.alanba.com', 'gradworks.umi.com', 'books.google.com', 'books.google.com', 'www.steelorbis.com', 'query.nytimes.com', 'theconversation.com', 'www.process-worldwide.com', 'books.google.com', 'www.usatoday.com', 'www.britannica.com', 'beltandroad.hktdc.com', 'gulfnews.com', 'www.constructionweekonline.com', 'www.bloomberg.com', 'books.google.com', 'encarta.msn.com', 'books.google.com', 'www.aljazeera.com', 'www.birdguides.com', 'books.google.com', 'news.satnews.com', 'www.alraimedia.com', 'www.youtube.com', 'www.al-monitor.com', 'www.spglobal.com', 'books.google.com', 'www.constructionweekonline.com', 'spacenews.com', 'www.thefreelibrary.com', 'www.nesfircroft.com', 'www.nytimes.com', 'www.constructionweekonline.com', 'www.unesco.org', 'rsf.org', 'www.jstor.org', 'www.imf.org', 'www.socialprogress.org', 'darmuseum.org', 'network.satnogs.org', 'freedomhouse.org', 'unpan1.un.org', 'www.washingtoninstitute.org', 'undocs.org', 'www.atlanticcouncil.org', 'data.footprintnetwork.org', 'www.unhcr.org', 'carnegieendowment.org', 'www.artkuwait.org', 'www.hrw.org', 'rsf.org', 'www.washingtoninstitute.org', 'services.tsck.org', 'www.un.org', 'data.worldbank.org', 'jstor.org', 'kfas.org', 'meetingorganizer.copernicus.org', 'www.hospitalitynet.org', 'www.amar-foundation.org', 'hdr.undp.org', 'widgets.weforum.org', 'hdr.undp.org', 'www.imf.org', 'www.transparency.org', 'www.imf.org', 'darmuseum.org', 'whc.unesco.org', 'nationalinterest.org', 'rsf.org', 'www.sesrtcic.org', 'www.freedomhouse.org', 'fpif.org', 'www.wttc.org', 'reports.weforum.org', 'fred.stlouisfed.org', 'en.unesco.org', 'darmuseum.org', 'www.orbitalspace.org', 'uprdoc.ohchr.org', 'www.ameu.org', 'hdr.undp.org', 'rsf.org', 'www.humanrightsfirst.org', 'babel.hathitrust.org', 'www.hrw.org', 'www.porttechnology.org', 'www.unesco.org', 'avibase.bsc-eoc.org', 'www.agsiw.org', 'www.archaeology.org', 'freedomhouse.org', 'www.systemicpeace.org', 'kfas.org', 'www.hrw.org', 'data.worldbank.org', 'ed-thelen.org', 'kottke.org', 'datazone.birdlife.org', 'www.constituteproject.org', 'globalsecurity.org', 'www.oxgaps.org', 'www.jstor.org', 'feow.org', 'www.ibe.unesco.org', 'darmuseum.org', 'www.refworld.org', 'www.archaeology.org', 'www.swfinstitute.org', 'www.amar-foundation.org', 'carnegieendowment.org', 'oxgaps.org', 'rsf.org', 'www.ibraaz.org', 'www.fao.org', 'www.unescwa.org', 'www.refworld.org', 'www.freedomhouse.org', 'warehouse.funcube.org', 'science.org', 'arteeast.org', 'freedomhouse.org', 'rsf.org', 'freedomhouse.org', 'www.fao.org', 'www.artpapers.org', 'freedomhouse.org', 'freedomhouse.org', 'en.wikisource.org', 'artkuwait.org', 'rsf.org', 'acig.org', 'www.artpapers.org', 'www.kfas.org', 'hdr.undp.org', 'survey07.ituc-csi.org', 'rsf.org', 'www.mcquaid.org', 'www.un.org', 'www.systemicpeace.org', 'www.aaa.org', ['[[bmc health services research'], ['archaeology international'], ['annals of clinical psychiatry'], ['quaternary research'], ['education as change'], ['arabian archaeology and epigraphy'], ['british journal of middle eastern studies'], ['built environment '], ['british journal of middle eastern studies'], ['contemporary review of the middle east'], [' arabian archaeology and epigraphy'], ['dyslexia'], ['resources'], ['[[comparative studies of south asia'], ['desalination'], ['middle eastern studies'], ['arabian archaeology and epigraphy'], ['aquatic ecosystem health '], ['all azimuth'], ['jacques connan']]",7515890,Allow all users (no expiry set),283280,11 May 2001,KoyaanisQatsi ,10786,90,2001-05-11,2001-05,2001
314,314,Berlin,https://en.wikipedia.org/wiki/Berlin,289,0,[],[],16,1,0,94,0,3,176,0.05536332179930796,0.0034602076124567475,0.32525951557093424,0.0,0.0,0.058823529411764705,0,"['ftp.atdd.noaa.gov', 'www.economist.com', 'washingtonpost.com', 'foodtank.com', 'luxeadventuretraveler.com', 'www.nytimes.com', 'travelinho.com', 'travel.nytimes.com', 'euractiv.com', 'www.weatherbase.com', 'www.decodedmagazine.com', 'www.bloomberg.com', 'www.dw.com', 'books.google.com', 'books.google.com', 'de.statista.com', 'embassypages.com', 'www.bostonglobe.com', 'www.deutschebahn.com', 'books.google.com', 'www.nytimes.com', 'www.observer.com', 'www.handelsblatt.com', 'www.metrotimes.com', 'www.businessinsider.com', 'www.dw.com', 'www.nytimes.com', 'books.google.com', 'travel2.nytimes.com', 'books.google.com', 'mobilityexchange.mercer.com', 'www.fifa.com', 'www.wsj.com', 'www.siemens.com', 'www.saveur.com', 'www.newsweek.com', 'books.google.com', 'edition.cnn.com', 'weather.com', 'www.kpmg.com', 'www.nbcnews.com', 'www.weather-atlas.com', 'www.nytimes.com', 'books.google.com', 'www.expatica.com', 'www.nytimes.com', 'scc-events.com', 'www.bbc.com', 'travel2.nytimes.com', 'www.berliner-extremwerte.com', 'www.thejewishweek.com', 'www.dw.com', 'monocle.com', 'www.western-allies-berlin.com', 'blogs.bettor.com', 'de.statista.com', 'www.weatherbase.com', 'www.nytimes.com', 'travel2.nytimes.com', 'books.google.com', 'guide.michelin.com', 'www.slowtravelberlin.com', 'www.treehugger.com', 'www.iccaworld.com', 'www.credit-suisse.com', 'global.handelsblatt.com', 'www.time.com', 'travel2.nytimes.com', 'www.forbes.com', 'bayer.com', 'monocle.com', 'www.nytimes.com', 'travel2.nytimes.com', 'www.businessweek.com', 'www.nytimes.com', 'russiajournal.com', 'www.observer.com', 'www.cnn.com', 'citymayors.com', 'www.nytimes.com', 'www.huffingtonpost.com', 'books.google.com', 'www.bbc.com', 'www.natureindex.com', 'www.hubculture.com', 'de.statista.com', 'www.google.com', 'www.theage.com', 'www.newyorker.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.nytimes.com', 'bloomberg.com', 'www.telecompaper.com', 'whc.unesco.org', 'whc.unesco.org', 'whc.unesco.org', 'wayback.archive-it.org', 'www.metropolis2005.org', 'hdi.globaldatalab.org', 'www.ushmm.org', 'www.germanfoods.org', 'berlin2009.org', 'www.specialolympics.org', 'www.europeanfilmacademy.org', 'www.worldcat.org', 'www.h-net.org', 'www.deutsche-metropolregionen.org', 'www.worldweather.org', 'www.metropolis2005.org']",3354,Allow all users (no expiry set),231991,11 November 2001,H. Jonat~enwiki ,13293,14,2001-11-11,2001-11,2001
315,315,Matera,https://en.wikipedia.org/wiki/Matera,26,0,[],[],1,0,0,10,0,0,15,0.038461538461538464,0.0,0.38461538461538464,0.0,0.0,0.038461538461538464,0,"['italianfoodexcellence.com', 'books.google.com', 'lalucana.com', 'patch.com', 'videostatic.com', 'materaprivatetours.com', 'books.google.com', 'made-in-italy.com', 'divento.com', 'books.google.com', 'www.wmf.org']",60040,Allow all users (no expiry set),28992,20 June 2002,Vincenzo~enwiki ,612,0,2002-06-20,2002-06,2002
316,316,Antakya,https://en.wikipedia.org/wiki/Antakya,18,0,[],[],0,0,0,12,0,0,6,0.0,0.0,0.6666666666666666,0.0,0.0,0.0,0,"['www.aljazeera.com', 'books.google.com', 'books.google.com', 'books.google.com', 'edgeofhumanity.com', 'www.weatherbase.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'biblehub.com']",394998,Allow all users (no expiry set),30184,9 December 2003,Adam Bishop ,724,0,2003-12-09,2003-12,2003
317,317,Monza,https://en.wikipedia.org/wiki/Monza,8,0,[],[],0,0,0,2,0,0,6,0.0,0.0,0.25,0.0,0.0,0.0,0,"['www.heraldscotland.com', 'enterf1.com']",65143,Allow all users (no expiry set),32677,25 March 2002,Dch ,790,3,2002-03-25,2002-03,2002
318,318,Chhattisgarh,https://en.wikipedia.org/wiki/Chhattisgarh,94,0,[],[],8,19,0,34,0,0,33,0.0851063829787234,0.20212765957446807,0.3617021276595745,0.0,0.0,0.2872340425531915,0,"['www.censusindia.gov', 'industries.cg.gov', 'censusindia.gov', 'bastar.gov', 'india-wris.nrsc.gov', 'chhattisgarhmines.gov', 'censusindia.gov', 'india.gov', 'durg.gov', 'www.censusindia.gov', 'durg.gov', 'censusindia.gov', 'cg.gov', 'kanker.gov', 'cg.gov', 'cg.gov', 'www.secr.indianrailways.gov', 'censusindia.gov', 'uidai.gov', 'www.naidunia.com', 'www.haribhoomi.com', 'www.patrika.com', 'mapsofindia.com', '36.gurturgoth.com', 'timesofindia.indiatimes.com', 'zeenews.india.com', 'www.thehindu.com', 'cgclimatechange.com', 'swachhindia.ndtv.com', 'economictimes.indiatimes.com', 'kosalkatha.com', 'www.mapsofindia.com', 'www.dailypioneer.com', 'www.dailypioneer.com', 'www.dailypioneer.com', 'zeenews.india.com', '36.gurturgoth.com', 'books.google.com', 'www.populationu.com', 'books.google.com', 'tribes-of-india.blogspot.com', 'www.maniactravellers.com', 'www.districtsofindia.com', '36.gurturgoth.com', 'www.korbacity.com', 'www.maniactravellers.com', 'languageinindia.com', 'www.business-standard.com', 'www.google.com', 'swachhindia.ndtv.com', 'www.mapsofindia.com', 'www.mapsofindia.com', 'naidunia.jagran.com', 'www.downtoearth.org', 'prsindia.org', 'headlinestoday.org', 'globaldatalab.org', 'indiawaterportal.org', 'www.prsindia.org', 'www.wisdomlib.org', 'www.sangeetnatak.org']",47734,Allow all users (no expiry set),98995,5 April 2002,194.65.14.70 ,4242,12,2002-04-05,2002-04,2002
319,319,Telangana,https://en.wikipedia.org/wiki/Telangana,132,4,"['10.1017/s0021911800154841', '10.2307/2753831', '10.2307/2052408', '10.1017/s0026749x00004996', None, None, None, None, None, None, None, None]","[['the journal of asian studies ', 'association for asian studies '], ['pacific affairs ', 'university of british columbia '], ['journal of asian studies '], ['[[cambridge university press', '[[modern asian studies']]",9,22,0,69,0,0,28,0.06818181818181818,0.16666666666666666,0.5227272727272727,0.030303030303030304,0.0,0.26515151515151514,4,"['www.telangana.gov', 'www.telangana.gov', 'censusindia.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'www.scr.indianrailways.gov', 'newdistrictsformation.telangana.gov', 'www.telangana.gov', 'www.aponline.gov', 'www.telangana.gov', 'www.telangana.gov', 'apind.gov', 'www.roadbuild.telangana.gov', 'www.aponline.gov', 'www.aponline.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'ecostat.telangana.gov', 'www.scr.indianrailways.gov', 'apsrtc.gov', 'pib.gov', 'telangana.gov', 'telanganatoday.com', 'www.hindu.com', 'timesofindia.indiatimes.com', 'indianexpress.com', 'books.google.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.dnaindia.com', 'www.rediff.com', 'www.newindianexpress.com', 'www.thehindu.com', 'www.languageinindia.com', 'books.google.com', 'www.hindu.com', 'timesofindia.indiatimes.com', 'www.hyderabadisearch.com', 'timesofindia.indiatimes.com', 'www.britannica.com', 'www.outlookindia.com', 'www.thehindu.com', 'www.thehindubusinessline.com', 'www.thehansindia.com', 'hindu.com', 'www.hindustantimes.com', 'scclmines.com', 'www.newindianexpress.com', 'www.newindianexpress.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'www.politicsdaily.com', 'www.thehindu.com', 'www.thehansindia.com', 'telangana.pscnotes.com', 'timesofindia.indiatimes.com', 'www.siasat.com', 'news.google.com', 'books.google.com', 'www.thehindubusinessline.com', 'www.newindianexpress.com', 'www.dnaindia.com', 'timesofindia.indiatimes.com', 'www.deccanchronicle.com', 'www.thehindubusinessline.com', 'indiansaga.com', 'indianexpress.com', 'www.ndtv.com', 'www.deccanchronicle.com', 'www.thehindu.com', 'www.thehindubusinessline.com', 'www.thehindu.com', 'articles.economictimes.indiatimes.com', 'telanganatoday.com', 'insideismailism.files.wordpress.com', 'www.hindu.com', 'guinnessworldrecords.com', 'mahabubnagar.tripod.com', 'www.business-standard.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'www.thenewsminute.com', 'www.news18.com', 'timesofindia.indiatimes.com', 'ndtv.com', 'www.thehansindia.com', 'www.telanganastateinfo.com', 'www.templenet.com', 'www.apsmfc.com', 'whc.unesco.org', 'swaminomics.org', 'whc.unesco.org', 'www.telanganalegislature.org', 'www.rbi.org', 'himalayanconnections.org', 'hdi.globaldatalab.org', 'www.metmuseum.org', 'indianheartassociation.org', ['the journal of asian studies ', 'association for asian studies '], ['pacific affairs ', 'university of british columbia '], ['journal of asian studies '], ['[[cambridge university press', '[[modern asian studies']]",990267,Allow all users (no expiry set),110244,16 September 2004,Tom Radulovich ,8704,12,2004-09-16,2004-09,2004
320,320,Jodhpur,https://en.wikipedia.org/wiki/Jodhpur,51,0,[],[],1,12,0,30,0,0,8,0.0196078431372549,0.23529411764705882,0.5882352941176471,0.0,0.0,0.2549019607843137,0,"['jda.urban.rajasthan.gov', 'urban.rajasthan.gov', 'jda.urban.rajasthan.gov', 'amssdelhi.gov', 'www.censusindia.gov', 'imdpune.gov', 'censusofindia.gov', 'jda.urban.rajasthan.gov', 'imdpune.gov', 'imdpune.gov', 'jda.urban.rajasthan.gov', 'jodhpur.rajasthan.gov', 'www.patrika.com', 'www.firstpost.com', 'www.patrika.com', 'books.google.com', 'www.nytimes.com', 'timesofindia.indiatimes.com', 'epaper.dainikjaltedeep.com', 'www.forbesindia.com', 'www.dnaindia.com', 'zeenews.india.com', 'books.google.com', 'www.timesofindia.com', 'indiarailinfo.com', 'www.outlookindia.com', 'www.thehindubusinessline.com', 'articles.timesofindia.indiatimes.com', 'www.amarujala.com', 'hindi.news18.com', 'www.dnaindia.com', 'www.bhaskar.com', 'www.timesofindia.com', 'www.bhaskar.com', 'www.huffpost.com', 'webconte.com', 'india.com', 'food.ndtv.com', 'indianexpress.com', 'www.bhaskar.com', 'www.bhaskar.com', 'www.indiatvnews.com', 'jodhpurmc.org']",983053,Allow all users (no expiry set),53245,13 September 2004,LeeHunter ,3311,6,2004-09-13,2004-09,2004
321,321,Bari,https://en.wikipedia.org/wiki/Bari,28,1,"['10.1080/00420988520080361', None, None]",[['urban studies ']],1,0,0,10,0,0,17,0.03571428571428571,0.0,0.35714285714285715,0.03571428571428571,0.0,0.07142857142857142,1,"['news.google.com', 'www.moovitapp.com', 'www.com', 'books.google.com', 'www.amazon.com', 'www.moovitapp.com', 'www.mapquest.com', 'www.com', 'www.com', 'www.britannica.com', 'creativecommons.org', ['urban studies ']]",44784,Allow all users (no expiry set),43023,18 March 2002,62.98.20.244 ,1294,1,2002-03-18,2002-03,2002
322,322,Haryana,https://en.wikipedia.org/wiki/Haryana,239,0,[],[],10,44,0,137,0,0,49,0.04184100418410042,0.18410041841004185,0.5732217573221757,0.0,0.0,0.22594142259414227,0,"['www.schooleducationharyana.gov', 'hpgcl.gov', 'censusindia.gov', 'imdpune.gov', 'dfccil.gov', 'www.nwr.indianrailways.gov', 'www.haryana.gov', 'haryanapoliceonline.gov', 'haryanatourism.gov', 'haryanatourism.gov', 'www.nr.indianrailways.gov', 'haryanaforest.gov', 'ncr.indianrailways.gov', 'csharyana.gov', 'hryedumis.gov', 'www.censusindia.gov', 'www.wii.gov', 'www.ncr.indianrailways.gov', 'haryanaforest.gov', 'dfccil.gov', 'www.schooleducationharyana.gov', 'india-wris.nrsc.gov', 'www.nr.indianrailways.gov', 'haryanacmoffice.gov', 'haryanatourism.gov', 'www.nr.indianrailways.gov', 'www.nwr.indianrailways.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'www.nrhm.gov', 'www.indianrailways.gov', 'www.schooleducationharyana.gov', 'www.cr.indianrailways.gov', 'www.indianrail.gov', 'censusindia.gov', 'www.nwr.indianrailways.gov', 'haryanaforest.gov', 'www.pmindia.gov', 'imdpune.gov', 'haryanaforest.gov', 'india.gov', 'www.haryanatourism.gov', 'haryanaforest.gov', 'www.haryana.gov', 'indianexpress.com', 'cities.expressindia.com', 'www.business-standard.com', 'www.hindustantimes.com', 'www.hindustantimes.com', 'www.hccinfrastructure.com', 'www.indiaclub.com', 'www.indianexpress.com', 'www.uniindia.com', 'indianexpress.com', 'www.tribuneindia.com', 'www.jagran.com', 'www.indianexpress.com', 'www.jagran.com', 'books.google.com', 'timesofindia.indiatimes.com', 'unemploymentinindia.cmie.com', 'books.google.com', 'indianexpress.com', 'books.google.com', 'indianexpress.com', '2fwww.jagran.com', 'cities.expressindia.com', 'www.travelbizmonitor.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.indianmirror.com', 'articles.economictimes.indiatimes.com', 'haryana-online.com', 'www.tribuneindia.com', 'content-www.cricinfo.com', 'domainmarket.com', 'haryana-online.com', 'books.google.com', 'haribhoomi.com', 'indianexpress.com', 'books.google.com', 'www.hindustantimes.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.thehindubusinessline.com', 'www.hillsofmorni.com', 'books.google.com', 'books.google.com', 'www.hindustantimes.com', 'in.jagran.yahoo.com', 'www.tribuneindia.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.dailypioneer.com', 'books.google.com', 'www.forbes.com', 'www.vedamsbooks.com', 'articles.economictimes.indiatimes.com', 'books.google.com', 'www.hindustantimes.com', 'books.google.com', 'indianexpress.com', 'www.vedamsbooks.com', 'articles.timesofindia.indiatimes.com', 'www.tribuneindia.com', 'content-www.cricinfo.com', 'timesofindia.indiatimes.com', 'www.indianexpress.com', 'www.havells.com', 'www.ethnologue.com', 'books.google.com', 'cities.expressindia.com', 'news.webindia123.com', 'www.tribuneindia.com', 'www.dailypioneer.com', 'www.tribuneindia.com', 'zeenews.india.com', 'india.com', 'www.hindustantimes.com', 'www.tribuneindia.com', 'www.hindustantimes.com', 'www.tribuneindia.com', 'atlascyclesonepat.com', 'www.indianexpress.com', 'www.osramindia.com', 'books.google.com', 'news.google.com', 'www.tribuneindia.com', 'books.google.com', 'timesofindia.indiatimes.com', 'pressreader.com', 'books.google.com', 'www.thehindu.com', 'www.business-standard.com', 'timesofindia.indiatimes.com', 'eceindustriesltd.com', 'www.ijrsr.com', 'www.knowmyindia.com', 'books.google.com', 'books.google.com', 'books.google.com', 'haryanasamanyagyan.com', 'epaper.timesofindia.com', 'www.tribuneindia.com', 'www.thehindu.com', 'archive.indianexpress.com', 'www.tribuneindia.com', 'www.tribuneindia.com', 'www.axonvet.com', 'haryana-online.com', 'articles.economictimes.indiatimes.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.hindustantimes.com', 'books.google.com', 'books.google.com', 'economictimes.indiatimes.com', 'books.google.com', 'hillsofmorni.com', 'www.haryana-online.com', 'books.google.com', 'books.google.com', 'iitd.ac.com', 'books.google.com', 'www.business-standard.com', 'www.dnaindia.com', 'www.damdamalake.com', 'books.google.com', 'lntgulf.com', 'www.tribuneindia.com', 'quickgs.com', 'books.google.com', 'www.indianexpress.com', 'www.hillsofmorni.com', 'books.google.com', 'timesofindia.indiatimes.com', 'punjabnewsline.com', 'books.google.com', 'cities.expressindia.com', 'www.ibef.org', 'www.isprs.org', 'www.downtoearth.org', 'wayback.archive-it.org', 'hdi.globaldatalab.org', 'www.icfa.org', 'www.bseh.org', 'www.isprs.org', 'www.haryanainvest.org', 'threatenedtaxa.org']",14189,Allow all users (no expiry set),156001,24 November 2001,Hagedis ,5609,34,2001-11-24,2001-11,2001
323,323,Sub-Saharan Africa,https://en.wikipedia.org/wiki/Sub-Saharan_Africa,256,15,"['10.1080/13629387.2011.635450', '10.1029/1999gl900494', '10.1016/j.tree.2018.05.005', '10.1126/science.aao6266', '10.1038/s41467-019-11213-w', '10.1038/194201a0', '10.3213/1612-1651-10153', '10.1126/science.1172257', '10.3213/1612-1651-10171', '10.1016/j.vaccine.2011.12.123', '10.1002/(sici)1099-1751(199706)12:1+<s29::aid-hpm465>3.0.co;2-u', '10.4135/9781452231648', '10.2307/1166258', '10.1080/13629387.2010.486573', '10.1086/505436', None, None, '30007846', '28971970', '31506422', None, None, '19407144', None, '22230581', '10173105', None, None, None, '16826514', None, None, '6092560', None, '6736881', None, None, '2947357', None, None, None, None, None, None, '1559480']","[['the journal of north african studies '], ['geophysical research letters '], ['trends in ecology '], ['science '], ['[[nature communications'], ['nature '], ['journal of african archaeology'], ['science '], ['[[journal of african archaeology'], ['vaccine '], ['the international journal of health planning and management '], ['sage publications'], ['issue'], ['the journal of north african studies '], ['the american journal of human genetics ']]",54,37,0,57,0,3,92,0.2109375,0.14453125,0.22265625,0.05859375,0.0,0.4140625,15,"['www.cia.gov', 'minerals.usgs.gov', 'www.csa.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'minerals.usgs.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.nigerianstat.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'minerals.usgs.gov', 'cia.gov', 'usaid.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'cia.gov', 'buanews.gov', 'minerals.usgs.gov', 'www.dst.gov', 'www.cia.gov', 'books.google.com', 'www.bbportuguese.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.sciencedaily.com', 'www.theatlantic.com', 'books.google.com', 'www.gallup.com', 'blogspot.com', 'www.sciencefriday.com', 'books.google.com', 'books.google.com', 'www.economist.com', 'sciencedaily.com', 'www.nytimes.com', 'site.ebrary.com', 'books.google.com', 'www.fasken.com', 'gold-eagle.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.ethnologue.com', 'www.nytimes.com', 'books.google.com', 'www.africannewsworld.com', 'allafrica.com', 'about.com', 'books.google.com', 'www.thelanguagejournal.com', 'books.google.com', 'www.economist.com', 'books.google.com', 'www.foreignpolicy.com', 'books.google.com', 'redorbit.com', 'www.sciencedaily.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.pulseafrica.com', 'www.nytimes.com', 'www.sportsscientists.com', 'upi.com', 'works.bepress.com', 'mbendi.com', 'books.google.com', 'worlddefensereview.com', 'books.google.com', 'killerplants.com', 'books.google.com', 'books.google.com', 'esa.un.org', 'data.worldbank.org', 'unaids.org', 'monthlyreview.org', 'unesdoc.unesco.org', 'www.unaids.org', 'world-nuclear.org', 'infosamak.org', 'iaaf.org', 'metmuseum.org', 'www.unaids.org', 'worldbank.org', 'www.unesco.org', 'en.unesco.org', 'www.transparency.org', 'www.eib.org', 'www.pewforum.org', 'www.odi.org', 'transparency.org', 'www.cgdev.org', 'www.metmuseum.org', 'unstats.un.org', 'www.africanrockart.org', 'www.pambazuka.org', 'www.africa.undp.org', 'www.eldis.org', 'www.saylor.org', 'unstats.un.org', 'www.doingbusiness.org', 'www.unesco.org', 'infosamak.org', 'www.desmondtutuhivcentre.org', 'esa.un.org', 'wayback.archive-it.org', 'cdcdevelopmentsolutions.org', 'unesdoc.unesco.org', 'www.unesco.org', 'iaaf.org', 'secid.org', 'monthlyreview.org', 'dictionary.cambridge.org', 'www.unaids.org', 'www.worldbank.org', 'data.worldbank.org', 'somraf.org', 'data.worldbank.org', 'www-wds.worldbank.org', 'www.pambazuka.org', 'ng.boell.org', 'www.iea.org', 'www.prb.org', 'data.worldbank.org', 'pewforum.org', 'worldbank.org', ['the journal of north african studies '], ['geophysical research letters '], ['trends in ecology '], ['science '], ['[[nature communications'], ['nature '], ['journal of african archaeology'], ['science '], ['[[journal of african archaeology'], ['vaccine '], ['the international journal of health planning and management '], ['sage publications'], ['issue'], ['the journal of north african studies '], ['the american journal of human genetics ']]",27067,Allow all users (no expiry set),211108,25 February 2002,Conversion script ,4229,3,2002-02-25,2002-02,2002
324,324,Culture of Bulgaria,https://en.wikipedia.org/wiki/Culture_of_Bulgaria,33,0,[],[],6,1,0,10,0,0,16,0.18181818181818182,0.030303030303030304,0.30303030303030304,0.0,0.0,0.21212121212121213,0,"['lcweb2.loc.gov', 'www.bulgariainside.com', 'www.dramavarna.com', 'slusham.com', 'www.ploshtadslaveikov.com', 'www.teatarvtarnovo.com', 'novinite.com', 'www.britannica.com', 'www.bg-istoria.com', 'grammy.com', 'books.google.com', 'www.forum18.org', 'www.soros.org', 'young-bulgarian-artists.org', 'www.arttoday.org', 'ica-sofia.org', 'shechen-bg.org']",251620,Allow all users (no expiry set),40819,23 June 2003,136.142.22.230 ,368,1,2003-06-23,2003-06,2003
325,325,Milan,https://en.wikipedia.org/wiki/Milan,237,0,[],[],11,3,0,68,0,0,155,0.046413502109704644,0.012658227848101266,0.2869198312236287,0.0,0.0,0.05907172995780591,0,"['earthobservatory.nasa.gov', 'www1.interno.gov', 'www.gov', 'www.italianbusinesstips.com', 'britannica.com', 'www.cronicajalisco.com', 'www.accuweather.com', 'www.com', 'www.britannica.com', 'books.google.com', 'www.collinsdictionary.com', 'mediagallery.com', 'www.hindustantimes.com', 'www.demographia.com', 'magazine.fourseasons.com', 'www.trenitalia.com', 'frieze.com', 'explo-re.com', 'www.languagemonitor.com', 'statista.com', 'mojeh.com', 'www.accuweather.com', '100milano.com', 'lankaramaya.com', 'euromonitor.com', 'www.forbes.com', 'www.com', 'www.bbc.com', 'archdaily.com', 'www.com', 'frogdesign.com', 'explo-re.com', 'www.statista.com', 'gamesbids.com', 'holyday-weather.com', 'unseendestination.com', 'www.com', 'rankings.ft.com', 'money.cnn.com', 'www.topuniversities.com', 'www.com', 'www.scmp.com', 'books.google.com', 'rankings.ft.com', 'www.collinsdictionary.com', 'www.com', 'newsroom.mastercard.com', 'monocle.com', 'www.forbes.com', 'www.gam-milano.com', 'www.topuniversities.com', 'books.google.com', 'www.cavalleriasanmaurizio.com', 'weather-and-climate.com', 'news.microsoft.com', 'www.euronews.com', 'weatherspark.com', 'timeshighereducation.com', 'www.firstpost.com', 'www.italian-design-academy.com', 'www.google.com', 'books.google.com', 'languagemonitor.com', 'assaeroporti.com', 'gamesbids.com', 'pasticceriacova.com', 'www.group.intesasanpaolo.com', 'www.viamichelin.com', 'www.railwaygazette.com', 'www.nytimes.com', 'www.battlefieldanomalies.com', 'assets.pewresearch.org', 'ctbuh.org', 'milan.citylisting.org', 'www.ersa.org', 'unipiams.org', 'cambridge.org', 'www.esfr.org', 'www.oecd-ilibrary.org', 'newadvent.org', 'www.ismu.org', 'world.nycsubway.org']",36511,"Require autoconfirmed or confirmed access (15:14, 13 June 2022)",177416,4 February 2002,Derek Ross ,8935,4,2002-02-04,2002-02,2002
326,326,New England,https://en.wikipedia.org/wiki/New_England,194,3,"['10.1080/09658416.2021.2000996', '10.1017/s0021875812000709', None, None, None, '22145497', None, None, None]","[['language awareness '], ['journal of american studies'], ['national vital statistics reports']]",37,35,0,72,0,0,47,0.19072164948453607,0.18041237113402062,0.3711340206185567,0.015463917525773196,0.0,0.3865979381443299,3,"['www.census.gov', 'www.bea.gov', 'www.govinfo.gov', 'tigerweb.geo.census.gov', 'www2.census.gov', 'factfinder.census.gov', 'www.eia.doe.gov', 'ct.gov', 'factfinder.census.gov', 'www.loc.gov', 'factfinder.census.gov', 'factfinder.census.gov', 'sanders.senate.gov', 'factfinder.census.gov', 'factfinder.census.gov', 'www.nps.gov', 'www.census.gov', 'www.nass.usda.gov', 'water.usgs.gov', 'www.bls.gov', 'factfinder.census.gov', 'www.buyusa.gov', 'www.nass.usda.gov', 'www.nps.gov', 'www.census.gov', 'webarchive.loc.gov', 'www.bls.gov', 'www.nass.usda.gov', 'www.eia.doe.gov', 'factfinder.census.gov', 'www.bea.gov', 'factfinder.census.gov', 'www.census.gov', 'www.census.gov', 'www.nass.usda.gov', 'www.vhist.com', 'www.nytimes.com', 'encarta.msn.com', 'books.google.com', 'boston.com', 'u-s-history.com', 'www.concordmonitor.com', 'slavenorth.com', 'www.bostonmagazine.com', 'nes.com', 'www.salon.com', 'books.google.com', 'www.gallup.com', 'www.cnn.com', 'dictionary.reference.com', 'www.pressherald.com', 'www.thesportsdish.com', 'books.google.com', 'www.politico.com', 'masslive.com', 'courant.com', 'www.houghtonmifflinbooks.com', 'boston.com', 'www.britannica.com', 'britannica.com', 'www.fodors.com', 'boston.cbslocal.com', 'books.google.com', 'boston.com', 'www.boston.com', 'usatodayhss.com', 'thedailyreview.com', 'boston.com', 'athlonsports.com', 'salemwitchtrialsmuseum.com', 'www.boston.com', 'eagletribune.com', 'glo-con.com', 'www.zyen.com', 'www.allamericanpatriots.com', 'www.midcoast.com', 'books.google.com', 'books.google.com', 'books.google.com', 'chicagotribune.com', 'books.google.com', 'eagletribune.com', 'books.google.com', 'www.masscandlepin.com', 'www.courant.com', 'books.google.com', 'query.nytimes.com', 'www.gallup.com', 'newengland.com', 'www.boston.com', 'www.beeradvocate.com', 'books.google.com', 'www.scribd.com', 'www.usatoday.com', 'boston.com', 'www.nytimes.com', 'www.thefreedictionary.com', 'traveltips.usatoday.com', 'www.visitrhodeisland.com', 'www.bostonmagazine.com', 'encarta.msn.com', 'books.google.com', 'wallethub.com', 'omaha.com', 'gallup.com', 'www.britannica.com', 'books.google.com', 'discovernewengland.org', 'spectator.org', 'rhodetour.org', 'www.colonialwarsct.org', 'geology.teacherfriendlyguide.org', 'rhodetour.org', 'geology.teacherfriendlyguide.org', '(sechistorical.org', 'www.rihs.org', 'bostonfed.org', 'www.ncsl.org', 'www.bos.frb.org', 'www.poetryfoundation.org', 'www.profootballresearchers.org', 'www.masshist.org', 'www.jstor.org', 'taxhistory.org', 'ilsr.org', 'www.abenakination.org', 'quahog.org', 'www.ctheritage.org', 'abenakination.org', 'www.fenwayparkwriters.org', 'www.discovernewengland.org', 'www.flowofhistory.org', 'www.mountwashington.org', 'oldfilm.org', 'www.mountwashington.org', 'www.discovernewengland.org', 'www.harbus.org', 'colonialwarsct.org', 'nationalhumanitiescenter.org', 'scboston.org', 'needhamhistory.org', 'www.commonwealmagazine.org', 'www.bostonredevelopmentauthority.org', 'www.bpl.org', ['language awareness '], ['journal of american studies'], ['national vital statistics reports']]",21531764,Require administrator access (no expiry set),166796,5 February 2003,Sfmontyo ,8342,5,2003-02-05,2003-02,2003
327,327,Naples,https://en.wikipedia.org/wiki/Naples,205,3,"['10.2307/2547529', '10.3280/cad2015-001003', '10.2307/990664', None, None, None, None, None, None]","[['international migration review '], ['cadmo'], ['journal of the society of architectural historians ', 'university of california press ']]",7,1,0,90,0,2,103,0.03414634146341464,0.004878048780487805,0.43902439024390244,0.014634146341463415,0.0,0.05365853658536585,3,"['www.protezionecivile.gov', 'naples.rome-in-italy.com', 'books.google.com', 'www.bloomberg.com', 'books.google.com', 'books.google.com', 'www.reuters.com', 'moovitapp.com', 'books.google.com', 'cucinet.com', 'chabadnapoli.com', 'www.questia.com', 'books.google.com', 'books.google.com', 'www.fornobravo.com', 'about.com', 'www.com', 'www.com', 'books.google.com', 'holidaycityflash.com', 'railway-technology.com', 'www.questia.com', 'skyteam.com', 'www.com', 'www.com', 'books.google.com', 'timelineindex.com', 'naplesldm.com', 'planetware.com', 'naplesldm.com', 'www.com', 'books.google.com', 'www.red-travel.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.apimages.com', 'books.google.com', 'virtualtourist.com', 'naples.rome-in-italy.com', 'books.google.com', 'travel.nytimes.com', 'finefretted.com', 'grandi-tenori.com', 'naplesherald.com', 'www.com', 'ilgiornaledellarte.com', 'books.google.com', 'demotix.com', 'pizzatoday.com', 'naplesldm.com', 'www.com', 'goeurope.com', 'moovitapp.com', 'portanapoli.com', 'www.worldportsource.com', 'napoli2000.com', 'books.google.com', 'raileurope.com', 'naplesldm.com', 'lagunaguitars.com', 'www.britannica.com', 'www.apimages.com', 'www.imdb.com', 'books.google.com', 'about.com', 'www.britannica.com', 'student.britannica.com', 'classicalmusic.about.com', 'ethnologue.com', 'splendoroftruth.com', 'napoliaffari.com', 'naplesmylove.com', 'italianfoodforever.com', 'bellaonline.com', 'euromonitor.com', 'books.google.com', 'whatsonwhen.com', 'www.imdb.com', 'www.ukmediacentre.pwc.com', 'onestopitaly.com', 'www.com', 'onwar.com', 'www.com', 'bartleby.com', 'naplesldm.com', 'books.google.com', 'www.historytoday.com', 'earlyromanticguiar.com', 'www.com', 'en.com', 'azerbaijans.com', 'oah.org', 'wmflabs.org', 'www.unhabitat.org', 'creativecommons.org', 'www.sangennaro.org', 'seatemperature.org', 'www.theparisreview.org', ['international migration review '], ['cadmo'], ['journal of the society of architectural historians ', 'university of california press ']]",55880,Allow all users (no expiry set),165263,12 December 2001,64.210.248.xxx ,5641,11,2001-12-12,2001-12,2001
328,328,Mithila (region),https://en.wikipedia.org/wiki/Mithila_(region),37,0,[],[],1,0,0,22,0,1,13,0.02702702702702703,0.0,0.5945945945945946,0.0,0.0,0.02702702702702703,0,"['books.google.com', 'books.google.com', 'ndtv.com', 'books.google.com', 'kathmandupost.com', 'books.google.com', 'www.business-standard.com', 'books.google.com', 'newindianexpress.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.newindianexpress.com', 'kathmandupost.ekantipur.com', 'books.google.com', 'books.google.com', 'ekantipur.com', 'books.google.com', 'www.seasonsindia.com', 'books.google.com', 'www.anubhuti-hindi.org']",15128951,Allow all users (no expiry set),28005,9 January 2008,Pravinjha ,1000,13,2008-01-09,2008-01,2008
329,329,Molise,https://en.wikipedia.org/wiki/Molise,13,0,[],[],2,0,0,1,0,0,10,0.15384615384615385,0.0,0.07692307692307693,0.0,0.0,0.15384615384615385,0,"['www.collinsdictionary.com', 'hdi.globaldatalab.org', 'abruzzomoliseheritagesociety.org']",79641,Allow all users (no expiry set),22414,2 September 2002,64.157.78.106 ,688,0,2002-09-02,2002-09,2002
330,330,Tirana,https://en.wikipedia.org/wiki/Tirana,184,5,"['10.1080/13600820802090512', '10.1080/02665433.2011.601610', '10.1127/0941-2948/2006/0130', '10.1016/j.cities.2010.02.002', '10.1017/s0068245400019043', None, None, None, None, None, None, None, None, None, None]","[['global society'], ['planning perspectives '], ['[[meteorologische zeitschrift'], ['cities '], ['the annual of the british school at athens', 'british school at athens']]",13,21,0,49,0,3,93,0.07065217391304347,0.11413043478260869,0.266304347826087,0.02717391304347826,0.0,0.21195652173913043,5,"['www.instatgis.gov', 'www.tirana.gov', 'www.instat.gov', 'www.instat.gov', 'www.ata.gov', 'www.instat.gov', 'arsimi.gov', 'planifikimi.gov', 'www.instat.gov', 'www.instat.gov', 'www.instatgis.gov', 'www.tirana.gov', 'ata.gov', 'www.instat.gov', 'ftp.atdd.noaa.gov', 'www.instat.gov', 'english.beijing.gov', 'www.instat.gov', 'tirana.gov', 'www.state.gov', 'www.qarkutirane.gov', 'www.world-gazetteer.com', 'books.google.com', 'www.tiranatimes.com', 'www.youtube.com', 'www.arabianbusiness.com', 'www.biography.com', 'www.myalbanianfood.com', 'books.google.com', 'currentresults.com', 'www.gazeta-shqip.com', 'mobike.com', 'books.google.com', 'www.archdaily.com', 'www.panorama.com', 'www.euronews.com', 'www.nytimes.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'telegrafi.com', 'www.dw.com', 'www.com', 'www.nytimes.com', 'english.albeu.com', 'currentresults.com', 'www.tiranatimes.com', 'www.forum-al.com', 'www.youtube.com', 'www.weather-atlas.com', 'ecovolis.com', 'www.com', 'books.google.com', 'seenews.com', 'edition.cnn.com', 'sportekspres.com', 'www.nytimes.com', 'english.albeu.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'www.ocnal.com', 'forum-al.com', 'www.vogue.com', 'english.albeu.com', 'www.dw.com', 'www.reuters.com', 'ijbcnet.com', 'www.dw.com', 'articles.latimes.com', 'aam.org', 'aftirana.org', 'www.ecat-tirana.org', 'osce.org', 'www.fes-tirana.org', 'www.eltis.org', 'agroweb.org', 'www.annalindhfoundation.org', 'meteo-climat-bzh.dyndns.org', 'kryegjyshataboterorebektashiane.org', 'www.osce.org', 'www.osce.org', 'www.youthforum.org', ['global society'], ['planning perspectives '], ['[[meteorologische zeitschrift'], ['cities '], ['the annual of the british school at athens', 'british school at athens']]",31075,Require administrator access (no expiry set),127661,4 November 2001,ChuckSmith ,4705,0,2001-11-04,2001-11,2001
331,331,Copenhagen,https://en.wikipedia.org/wiki/Copenhagen,311,0,[],[],6,1,0,101,0,1,202,0.01929260450160772,0.003215434083601286,0.3247588424437299,0.0,0.0,0.022508038585209004,0,"['beijing.gov', 'books.google.com', 'www.tyznik.com', 'www.citymayors.com', 'danishnet.com', 'www.visitcopenhagen.com', 'www.visitcopenhagen.com', 'www.10kswim.com', 'www.visitcopenhagen.com', 'books.google.com', 'www.aljazeera.com', 'www.scandinaviastandard.com', 'www.moodiereport.com', 'travel.usnews.com', 'www.visitcopenhagen.com', 'www.cnn.com', 'www.railjournal.com', 'www.copcap.com', 'www.bbc.com', 'www.topuniversities.com', 'virgin-vacations.com', 'annualreport2012.cmport.com', 'books.google.com', 'www.architecture-page.com', 'www.shanghairanking.com', 'books.google.com', 'dualcitizeninc.com', 'finestclubs.com', 'www.copcap.com', 'www.topuniversities.com', 'www.nysun.com', 'www.welcome-to-my-copenhagen.com', 'books.google.com', 'britishbattles.com', 'www.carlsberggroup.com', 'dailyhomelist.com', 'arcspace.com', 'www.topuniversities.com', 'books.google.com', 'copenhagenfashionweek.com', 'books.google.com', 'flightstats.com', 'www.meetincopenhagen.com', 'www.weather-and-climate.com', 'books.google.com', 'www.forbes.com', 'emporis.com', 'www.visitcopenhagen.com', 'www.citymayors.com', 'www.visitcopenhagen.com', 'books.google.com', 'www.dezeen.com', 'books.google.com', 'arup.com', 'www.visitdenmark.com', 'books.google.com', 'visitcopenhagen.com', 'www.citymayors.com', 'books.google.com', 'www.visitcopenhagen.com', 'www.visitcopenhagen.com', 'www.neweuropeaneconomy.com', 'books.google.com', 'www.damvad.com', 'books.google.com', 'www.usatoday.com', 'books.google.com', 'books.google.com', 'www.visitcopenhagen.com', 'www.uefa.com', 'visitcopenhagen.com', 'www.travtasy.com', 'www.visitcopenhagen.com', 'books.google.com', 'books.google.com', 'voiceofrussia.com', 'railwaytechnology.com', 'www.henninglarsen.com', 'www.visitcopenhagen.com', 'books.google.com', 'worldhotels.com', 'www.henninglarsen.com', 'www.visitcopenhagen.com', 'books.google.com', 'www.nytimes.com', 'stateofgreen.com', 'www.visitcopenhagen.com', 'www.weather-atlas.com', 'www.visitcopenhagen.com', 'www.visitcopenhagen.com', 'danishnet.com', 'www.visitcopenhagen.com', 'books.google.com', 'www.visitcopenhagen.com', 'www.visitcopenhagen.com', 'books.google.com', 'books.google.com', 'www.visitdenmark.com', 'books.google.com', 'books.google.com', 'monocle.com', 'www.dictionary.com', 'www.oresundsregionen.org', 'meteo-climat-bzh.dyndns.org', 'www.opensocietyfoundations.org', 'dbs.bh.org', 'www.svoem.org', 'pub.nordregio.org']",5166,Require administrator access (no expiry set),228860,25 September 2001,194.95.63.xxx ,7679,5,2001-09-25,2001-09,2001
332,332,Königsberg,https://en.wikipedia.org/wiki/K%C3%B6nigsberg,132,1,"['10.1080/14650040903486967', None, None]",[['geopolitics']],3,0,0,8,0,0,120,0.022727272727272728,0.0,0.06060606060606061,0.007575757575757576,0.0,0.030303030303030304,1,"['books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.dw.com', 'visitkaliningrad.com', 'books.google.com', 'books.google.com', 'www.memorialmuseums.org', 'ibiblio.org', 'www.wilsoncenter.org', ['geopolitics']]",15413504,Allow all users (no expiry set),73608,30 July 2005,Laur ,1247,14,2005-07-30,2005-07,2005
333,333,Culture of Sri Lanka,https://en.wikipedia.org/wiki/Culture_of_Sri_Lanka,20,0,[],[],2,2,0,9,0,0,7,0.1,0.1,0.45,0.0,0.0,0.2,0,"['www.statistics.gov', 'www.cia.gov', 'gallup.com', 'books.google.com', 'books.google.com', 'www.infolanka.com', 'bookonsrilanka.files.wordpress.com', 'books.google.com', 'lankalibrary.com', 'lanka.com', 'books.google.com', 'mahavamsa.org', 'www.jstor.org']",3008201,Allow all users (no expiry set),31903,27 October 2005,64.231.195.228 ,736,1,2005-10-27,2005-10,2005
334,334,Culture of Italy,https://en.wikipedia.org/wiki/Culture_of_Italy,110,1,[],[],8,3,0,60,0,0,39,0.07272727272727272,0.02727272727272727,0.5454545454545454,0.00909090909090909,0.0,0.10909090909090909,0,"['state.gov', 'cia.gov', 'thomas.loc.gov', 'www.everyculture.com', 'unrv.com', 'books.google.com', 'scholastic.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.sorrisi.com', 'books.google.com', 'dot.com', 'books.google.com', 'wiley.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'www.topuniversities.com', 'books.google.com', 'books.google.com', 'frieze.com', 'books.google.com', 'scholastic.com', 'books.google.com', 'formula1.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.spainexchange.com', 'books.google.com', 'books.google.com', 'filmreference.com', 'shanghairanking.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'italoamericano.com', 'books.google.com', 'books.google.com', 'italytravel.com', 'www.spainexchange.com', 'books.google.com', 'topics.nytimes.com', 'books.google.com', 'books.google.com', 'cwur.org', 'whc.unesco.org', 'immaculateheartacademy.org', 'faostat.fao.org', 'faostat.fao.org', 'www.justitaly.org', 'pewforum.org', 'www.eoearth.org']",283846,Allow all users (no expiry set),140039,29 July 2003,Theanthrope ,4855,2,2003-07-29,2003-07,2003
335,335,Tourism in Lebanon,https://en.wikipedia.org/wiki/Tourism_in_Lebanon,47,1,"['10.1080/0966369x.2012.753586', None, None]",[['gender']],10,9,0,23,0,0,4,0.2127659574468085,0.19148936170212766,0.48936170212765956,0.02127659574468085,0.0,0.425531914893617,1,"['www.cas.gov', 'www.gov', 'www.destinationlebanon.gov', 'www.destinationlebanon.gov', 'travel.state.gov', 'www.destinationlebanon.gov', 'www.destinationlebanon.gov', 'www.destinationlebanon.gov', 'www.destinationlebanon.gov', 'www.mea.com', 'www.everyculture.com', 'about.com', 'www.forbes.com', 'www.travel-to-lebanon.com', 'lebanon.com', 'www.lebanonatlas.com', 'www.ikamalebanon.com', 'www.lebaneseexaminer.com', 'www.orient-latin.com', 'www.usatoday.com', 'www.travel-to-lebanon.com', 'orchid-lifestyle.com', 'www.rjliban.com', 'brite.blominvestbank.com', 'www.middleeast.com', 'www.travel-to-lebanon.com', 'www.nationsencyclopedia.com', 'www.soundcloud.com', 'a1-images.myspacecdn.com', 'www.menafn.com', 'www.sallys-place.com', 'abcnews.go.com', 'www.lebanonembassyus.org', 'whc.unesco.org', 'whc.unesco.org', 'whc.unesco.org', 'unwto.org', 'www.city-journal.org', 'whc.unesco.org', 'whc.unesco.org', 'unwto.org', 'whc.unesco.org', ['gender']]",13939289,Allow all users (no expiry set),79112,27 October 2007,Modar1hazar ,450,2,2007-10-27,2007-10,2007
336,336,Rum,https://en.wikipedia.org/wiki/Rum,76,1,"['10.1007/978-1-4615-0187-9_12', None, None]",[['springer']],2,1,0,17,0,0,55,0.02631578947368421,0.013157894736842105,0.2236842105263158,0.013157894736842105,0.0,0.05263157894736842,1,"['webarchive.nationalarchives.gov', 'www.scmp.com', 'liquor.com', 'www.oed.com', 'www.thrillist.com', 'www.westindiesrum.com', 'www.wired.com', '2fwww.snopes.com', 'www.bbc.com', 'books.google.com', 'www.hindu.com', 'the-rum-guys.com', 'blog.oup.com', 'www.oed.com', 'specialsections.nypost.com', 'www.sfgate.com', 'www.cigaraficionado.com', 'www.winemag.com', 'uniboa.org', 'www.fao.org', ['springer']]",14834691,Allow all users (no expiry set),47209,30 October 2001,212.248.133.xxx ,2540,7,2001-10-30,2001-10,2001
337,337,Bhutan,https://en.wikipedia.org/wiki/Bhutan,267,15,"['10.1080/13510347.2014.959437', '10.1017/s0030605300023619', '10.1093/jrs/9.4.397', '10.1038/s41467-020-19493-3', 'org/10.1093/jrs/9.4.397', '10.1057/9781137551429_1', '10.1111/j.1931-0846.2006.tb00521.x', '10.5502/ijw.v5i2.2', '10.1108/17465681211237600', '10.3390/resources7030058', '10.1080/0958493042000242954', '10.1108/gkmc-12-2019-0153', '10.1007/s10531-009-9587-5', '10.1896/052.023.0107', '10.1017/s0030605300033834', None, None, None, '33293507', None, None, None, None, None, None, None, None, None, None, None, None, None, None, '7723057', None, None, None, None, None, None, None, None, None, None, None]","[['democratization '], [' oryx '], ['journal of refugee studies '], ['nature communications'], ['journal of refugee studies'], ['palgrave macmillan'], ['geographical review '], ['international journal of wellbeing '], ['society and business review '], ['resources'], [' contemporary south asia '], ['global knowledge'], [' biodivers. conserv. '], [' primate conservation '], [' oryx ']]",59,19,0,108,0,3,64,0.2209737827715356,0.07116104868913857,0.4044943820224719,0.056179775280898875,0.0,0.34831460674157305,15,"['2001-2009.state.gov', 'www.mfa.gov', '2009-2017.state.gov', 'www.tourism.gov', 'www.gnhc.gov', 'www.acf.hhs.gov', 'www.cia.gov', 'www.westbengaltourism.gov', 'www.nab.gov', 'travel.state.gov', 'www.loc.gov', 'www.rcsc.gov', '2009-2017.state.gov', 'www.mfa.gov', 'www.loc.gov', 'www.bhutan.gov', 'state.gov', 'www.mfa.gov', '2001-2009.state.gov', 'books.google.com', 'books.google.com', 'www.climatechangenews.com', 'abroad.com', 'www.seattletimes.com', 'books.google.com', 'books.google.com', 'www.kuenselonline.com', 'www.bhutannewsservice.com', 'books.google.com', 'www.kuenselonline.com', 'www.kuenselonline.com', 'www.ambotravels.com', 'books.google.com', 'www.dhakatribune.com', 'www.ndtv.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.tribuneindia.com', 'www.dailybhutan.com', 'books.google.com', 'screamer.deadspin.com', 'books.google.com', 'www.seattletimes.com', 'www.atimes.com', 'www.cnn.com', 'www.techinasia.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'bdnews24.com', 'books.google.com', 'books.google.com', 'news.china.com', 'kuenselonline.com', 'www.holidify.com', 'www.scribd.com', 'www.ttgmice.com', 'www.britannica.com', 'books.google.com', 'en.prothom-alo.com', 'encarta.msn.com', 'www.impressbhutan.com', 'www.nytimes.com', 'bbc.com', 'books.google.com', 'www.dhakatribune.com', 'www.kuenselonline.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.bhutannewsservice.com', 'www.kuenselonline.com', 'www.nytimes.com', 'books.google.com', 'www.cnn.com', 'bhutantraveloperator.com', 'marktheday.com', 'www.tribuneindia.com', 'economictimes.indiatimes.com', 'books.google.com', 'www.digitalhimalaya.com', 'books.google.com', 'imnepal.com', 'ndtv.com', 'www.kuenselonline.com', 'www.kuenselonline.com', 'books.google.com', 'www.hindustantimes.com', 'www.kuenselonline.com', 'theweek.myrepublica.com', 'ngm.nationalgeographic.com', 'www.keystobhutan.com', 'www.kuenselonline.com', 'books.google.com', 'books.google.com', 'www.kuenselonline.com', 'www.gtpalliance.com', 'www.kuenselonline.com', 'books.google.com', 'www.upiasia.com', 'www.haaretz.com', 'timesofindia.indiatimes.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.bangkokpost.com', 'www.grossnationalhappiness.com', 'books.google.com', 'www.atimes.com', 'books.google.com', 'www.tribuneindia.com', 'www.oclarim.com', 'kuenselonline.com', 'www.ted.com', 'www.dnaindia.com', 'www.thimphutechpark.com', 'books.google.com', 'books.google.com', 'books.google.com', 'whc.unesco.org', 'www.wto.org', 'www.pri.org', 'www.adb.org', 'www.hydropower.org', 'www.unhcr.org', 'www.thlib.org', 'data.footprintnetwork.org', 'data.worldbank.org', 'www.pbs.org', 'www.worldinstituteforasianstudies.org', 'population.un.org', 'www.tradeforum.org', 'devdata.worldbank.org', 'data.worldbank.org', 'www.undp.org', 'www.worldwatchmonitor.org', 'hrw.org', 'asiasociety.org', 'whc.unesco.org', 'www.constituteproject.org', 'freedomhouse.org', 'www.hrw.org', 'www.amnesty.org', 'orientalbirdclub.org', 'www.imf.org', 'www.election-bhutan.org', 'whc.unesco.org', 'whc.unesco.org', 'minorityrights.org', 'sdfsec.org', 'www.refworld.org', 'hrw.org', 'whc.unesco.org', 'whc.unesco.org', 'www.amnesty.org', 'www.hrw.org', 'wdi.worldbank.org', 'whc.unesco.org', 'www.thlib.org', 'esa.un.org', 'hdr.undp.org', 'whc.unesco.org', 'esa.un.org', 'wdi.worldbank.org', 'www.bhutanstudies.org', 'hrw.org', 'www.bt.undp.org', 'www.thlib.org', 'www.un.org', 'www.hrw.org', 'esa.un.org', 'blogs.worldbank.org', 'www.democracy-international.org', 'www.adaptation-undp.org', 'www.unesco.org', 'www.pewforum.org', 'www.iucn.org', 'www.amnesty.org', ['democratization '], [' oryx '], ['journal of refugee studies '], ['nature communications'], ['journal of refugee studies'], ['palgrave macmillan'], ['geographical review '], ['international journal of wellbeing '], ['society and business review '], ['resources'], [' contemporary south asia '], ['global knowledge'], [' biodivers. conserv. '], [' primate conservation '], [' oryx ']]",2421391,Require administrator access (no expiry set),185016,22 April 2001,Koyaanisqatsi ,7027,44,2001-04-22,2001-04,2001
338,338,Indo-Persian culture,https://en.wikipedia.org/wiki/Indo-Persian_culture,17,0,[],[],4,0,0,3,0,0,10,0.23529411764705882,0.0,0.17647058823529413,0.0,0.0,0.23529411764705882,0,"['books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.iranicaonline.org', 'www.iranicaonline.org', 'www.iranicaonline.org', 'www.iranicaonline.org']",1291560,Allow all users (no expiry set),20249,17 December 2004,Sam Spade ,303,1,2004-12-17,2004-12,2004
339,339,Kannada people,https://en.wikipedia.org/wiki/Kannada_people,124,0,[],[],8,9,0,53,0,0,54,0.06451612903225806,0.07258064516129033,0.4274193548387097,0.0,0.0,0.13709677419354838,0,"['www.aponline.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'india.gov', 'ksdl.karnataka.gov', 'www.aponline.gov', 'www.censusindia.gov', 'censusindia.gov', 'archive.india.gov', 'www.rediff.com', 'timesofindia.indiatimes.com', 'books.google.com', 'archive.deccanherald.com', 'rediff.com', 'indiaprofile.com', 'timesofindia.indiatimes.com', 'www.hinduonnet.com', 'www.telegraphindia.com', 'www.hindu.com', 'daijiworld.com', 'archive.deccanherald.com', 'www.hindu.com', 'archive.deccanherald.com', 'www.ourkarnataka.com', 'pbs.twimg.com', 'www.caswath.com', 'www.gswift.com', 'archive.deccanherald.com', 'articles.timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.hindu.com', 'karnatakasanghamumbai.com', 'hindu.com', 'www.deccanherald.com', 'books.google.com', 'www.telegraphindia.com', 'temples.south-india-tour-package.com', 'lingayatreligion.com', 'www.templenet.com', 'atimes.com', 'www.kamat.com', 'hinduonnet.com', 'books.google.com', 'articles.timesofindia.indiatimes.com', 'www.deccanherald.com', 'www.lexico.com', 'www.pustakshakti.com', 'articles.timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.hindu.com', 'thehindu.com', 'books.google.com', 'www.ourkarnataka.com', 'encyclopedia.com', 'khadifederation.com', 'www.thehindu.com', 'www.deccanherald.com', 'www.hindu.com', 'newindianexpress.com', 'www.deccanchronicle.com', 'books.google.com', 'archive.deccanherald.com', 'www.kuwaitkannadakoota.org', 'singara.org', 'www.akkaonline.org', 'dallas.navika.org', 'sackannadasangha.org', 'www.nriforumkarnataka.org', 'www.singara.org', 'whc.unesco.org']",338799,Allow all users (no expiry set),69557,11 October 2003,Martalli ,2524,0,2003-10-11,2003-10,2003
340,340,Macedonians (ethnic group),https://en.wikipedia.org/wiki/Macedonians_(ethnic_group),245,18,"['10.1038/ejhg.2017.18', '10.1016/j.cub.2008.07.049', '10.1016/j.forsciint.2004.04.067', '10.1038/sj.ejhg.5200992', '10.1007/s10038-007-0125-6', '10.1038/ejhg.2014.50', '10.1371/journal.pone.0135820', '10.1111/j.1399-0039.2004.00273.x', '10.1038/nature07331', '10.1016/j.fsigen.2011.04.005', '10.15378/1848-9540.2014', '10.1080/0090599042000246406', '10.1163/187633004x00134', '10.1093/molbev/msi185', '10.1034/j.1399-0039.2000.550109.x', '10.1371/journal.pbio.1001555', '10.1126/science.290.5494.1155', None, '18691889', '15607593', '12825075', '17364156', '24667786', '26332464', '15361127', '18758442', '21549657', None, None, None, '15944443', '10703609', '23667324', '11073453', None, None, None, None, None, '4266736', '4558026', None, '2735096', None, None, None, None, None, None, '3646727', None]","[['[[european journal of human genetics'], ['curr. biol. '], [' forensic science international '], ['european journal of human genetics '], ['journal of human genetics'], [' european journal of human genetics '], [' plos one '], ['tissue antigens '], ['nature'], [' forensic sci. int. genet. '], [' etnološka tribina '], ['[[nationalities papers'], ['east central europe '], [' molecular biology and evolution '], ['tissue antigens'], ['[[plos biology'], ['science ']]",13,13,0,36,0,0,165,0.053061224489795916,0.053061224489795916,0.1469387755102041,0.07346938775510205,0.0,0.17959183673469387,17,"['www.censusdata.abs.gov', 'www.stats.gov', 'www.mfa.gov', 'www.mfa.gov', 'www.stat.gov', 'www.border.gov', 'www.census.gov', 'pod2.stat.gov', '2001-2009.state.gov', 'www.mfa.gov', 'www.mfa.gov', 'popis2021.stat.gov', 'www.census.gov', 'www.mia.com', 'balkaninsight.com', 'theconversation.com', 'www.kroraina.com', 'www.vreme.com', 'www.a1.com', 'books.google.com', 'books.google.com', 'www.dw.com', 'nationalpost.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.kroraina.com', 'www.etymonline.com', 'books.google.com', 'www.novamakedonija.com', 'www.utrinski.com', 'books.google.com', 'www.ethnologue.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.findarticles.com', 'books.google.com', 'www.findarticles.com', 'books.google.com', 'books.google.com', 'www.bbc.com', 'www.google.com', 'www.kroraina.com', 'books.google.com', 'books.google.com', 'gct.com', 'www.nytimes.com', 'www.monstat.org', 'www.amnesty.org', 'gbe.oxfordjournals.org', 'research.policyarchive.org', 'research.policyarchive.org', 'www.promacedonia.org', 'haemus.org', 'oscars.org', 'faq.macedonia.org', 'www.oecd.org', 'research.policyarchive.org', 'un.org', 'minorityrights.org', ['[[european journal of human genetics'], ['curr. biol. '], [' forensic science international '], ['european journal of human genetics '], ['journal of human genetics'], [' european journal of human genetics '], [' plos one '], ['tissue antigens '], ['nature'], [' forensic sci. int. genet. '], [' etnološka tribina '], ['[[nationalities papers'], ['east central europe '], [' molecular biology and evolution '], ['tissue antigens'], ['[[plos biology'], ['science ']]",432709,Require administrator access (no expiry set),137094,16 January 2004,217.79.65.243 ,7505,19,2004-01-16,2004-01,2004
341,341,Culture of the United Arab Emirates,https://en.wikipedia.org/wiki/Culture_of_the_United_Arab_Emirates,59,0,[],[],7,2,0,32,0,0,18,0.11864406779661017,0.03389830508474576,0.5423728813559322,0.0,0.0,0.15254237288135594,0,"['uae.gov', '2001-2009.state.gov', 'www.holidify.com', 'www.gulfnews.com', 'www.bayut.com', 'indexuae.com', 'gulfnews.com', 'gulfnews.com', 'www.commisceo-global.com', 'medium.com', 'www.bayut.com', 'books.google.com', 'uk.practicallaw.thomsonreuters.com', 'www.thenationalnews.com', 'www.commisceo-global.com', 'www.visitdubai.com', 'theculturetrip.com', 'books.google.com', 'uaeinteract.com', 'www.britannica.com', 'books.google.com', 'www.khaleejtimes.com', 'www.uaemoments.com', 'www.internationalcuisine.com', 'theculturetrip.com', 'www.thenationalnews.com', 'gulfnews.com', 'books.google.com', 'grapeshisha.com', 'www.yumpu.com', 'www.deezer.com', 'books.google.com', '200worldalbums.com', 'www.visitdubai.com', 'www.worldcat.org', 'archive.archaeology.org', 'www.uae-embassy.org', 'www.shayaan.org', 'www.worldcat.org', 'worldcat.org', 'earthsky.org']",20270829,Allow all users (no expiry set),28026,18 November 2008,TeamEnglish100Haven ,889,8,2008-11-18,2008-11,2008
342,342,Sinhalese people,https://en.wikipedia.org/wiki/Sinhalese_people,77,8,"[None, '10.1038/jhg.2013.112', '10.1002/ajpa.1330450112', '10.1086/499411', '10.1017/s0010417500017710', '10.1111/j.1744-313x.2007.00698.x', '10.2183/pjab.85.69', '10.1086/346068', '8908803', '24196378', None, '16400607', None, '17845299', '19212099', '12536373', None, None, None, '1380230', None, None, '3524296', '379225']","[['human biology '], ['journal of human genetics'], ['american journal of physical anthropology '], ['american journal of human genetics '], ['comparative studies in society and history'], ['international journal of immunogenetics '], ['proceedings of the japan academy. series b'], ['american journal of human genetics ']]",11,11,0,21,0,0,26,0.14285714285714285,0.14285714285714285,0.2727272727272727,0.1038961038961039,0.0,0.38961038961038963,8,"['www.statistics.gov', 'www.statistics.gov', 'www.stats.gov', 'www.statistics.gov', 'www.stats.gov', 'www.homeaffairs.gov', 'www.stats.gov', 'www.statistics.gov', 'www.dhs.gov', 'www.teara.gov', 'www.loc.gov', 'www.everyculture.com', 'www.lankalibrary.com', 'scenicsrilanka.com', 'lankalibrary.com', 'www.gallup.com', 'books.google.com', 'palikanon.com', 'sltouristguide.com', 'thestar.com', 'starofmysore.com', 'books.google.com', 'www.ethnologue.com', 'books.google.com', 'books.google.com', 'books.google.com', 'srilankanamericans.com', 'www.ethnologue.com', 'lankaemb-egypt.com', 'books.google.com', 'www.britannica.com', 's-media-cache-ak0.pinimg.com', 'mahavamsa.org', 'www.jstor.org', 'www.buddhistethics.org', 'www.jstor.org', 'isogg.org', 'mahavamsa.org', 'www.jstor.org', 'lakdiva.org', 'mahavamsa.org', 'angampora.org', 'www.kataragama.org', ['human biology '], ['journal of human genetics'], ['american journal of physical anthropology '], ['american journal of human genetics '], ['comparative studies in society and history'], ['international journal of immunogenetics '], ['proceedings of the japan academy. series b'], ['american journal of human genetics ']]",29359,Allow all users (no expiry set),59626,25 December 2001,213.17.74.xxx ,3259,3,2001-12-25,2001-12,2001
343,343,Gavar,https://en.wikipedia.org/wiki/Gavar,13,0,[],[],2,0,0,3,0,0,8,0.15384615384615385,0.0,0.23076923076923078,0.0,0.0,0.15384615384615385,0,"['www.findarmenia.com', 'www.kyavar.com', 'www.findarmenia.com', 'meteo-climat-bzh.dyndns.org', 'meteo-climat-bzh.dyndns.org']",2697674,Allow all users (no expiry set),20592,17 September 2005,24.205.21.196 ,305,0,2005-09-17,2005-09,2005
344,344,Somalis,https://en.wikipedia.org/wiki/Somalis,260,16,"['10.1371/journal.pgen.1004393', '10.1038/nature19310', '10.1086/382286', '10.1093/molbev/msm049', '10.1038/s41598-019-55344-y', '10.1007/978-90-481-2719-1_6', '10.1186/1471-2164-8-223', '10.1086/386294', '10.1038/ejhg.2008.70', '10.1038/s41598-020-62645-0', '10.3406/ethio.1976.1157', '10.1016/j.fsigen.2016.12.015', '10.1002/ajpa.20876', '10.1046/j.1529-8817.2003.00057.x', '10.1007/bf01540131', '10.1038/sj.ejhg.5201390', '24921250', '27459054', '14973781', '17351267', '31827175', None, '17620140', '15042509', '18398433', '32221414', None, '28068531', '18618658', '14748828', None, '15756297', '4055572', '5003663', '1182266', None, '6906521', None, '1945034', '1181964', None, '7101338', None, None, None, None, None, None]","[['plos genetics'], ['nature'], [' american journal of human genetics '], ['molecular biology and evolution'], ['scientific reports '], ['springer'], [' bmc genomics '], ['the american journal of human genetics'], ['european journal of human genetics '], ['scientific reports'], ['annales d'], ['forensic science international'], ['american journal of physical anthropology'], ['annals of human genetics '], ['computers and translation'], ['european journal of human genetics']]",19,9,0,73,0,0,144,0.07307692307692308,0.03461538461538462,0.28076923076923077,0.06153846153846154,0.0,0.16923076923076924,16,"['www.cia.gov', 'www.cia.gov', 'www.csa.gov', 'paperspast.natlib.gov', 'www.cia.gov', 'stats.gov', 'www.cia.gov', 'paperspast.natlib.gov', 'www.abs.gov', 'www.google.com', 'books.google.com', 'www.google.com', 'books.google.com', 'www.google.com', 'books.google.com', 'allafrica.com', 'www.ethnologue.com', 'www.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.nature.com', 'books.google.com', 'books.google.com', 'www.ethnologue.com', 'www.newspapers.com', 'lusakatimes.com', 'www.google.com', 'books.google.com', 'www.krepublishers.com', 'books.google.com', 'www.britannica.com', 'de.statista.com', 'www.google.com', 'www.citypages.com', 'ethnologue.com', 'books.google.com', 'www.docstoc.com', 'www.google.com', 'www.crwflags.com', 'www.independent.com', 'books.google.com', 'books.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.yfull.com', 'www.innercitypress.com', 'books.google.com', 'www.google.com', 'www.google.com', 'buluugleey.com', 'books.google.com', 'www.hiiraan.com', 'www.google.com', 'books.google.com', 'somalilandchronicle.com', 'books.google.com', 'www.ethnologue.com', 'foreignpolicy.com', 'www.fiba.com', 'books.google.com', 'www.google.com', 'www.google.com', 'books.google.com', 'books.google.com', 'jang.com', 'books.google.com', 'www.newspapers.com', 'www.hiiraan.com', 'www.omniglot.com', 'books.google.com', 'hiiraan.com', 'www.angelfire.com', 'books.google.com', 'strategypage.com', 'www.dawn.com', 'www.banadir.com', 'www.ethnologue.com', 'books.google.com', 'www.worldatlas.com', 'censusreporter.org', 'somalia.unfpa.org', 'karin-ha.org', 'www.un.org', 'www.un.org', 'www.hdcentre.org', 'unhcr.org', 'www.somaliweyn.org', 'peoplegroups.org', 'www.pewresearch.org', 'unhcr.org', 'peoplegroups.org', 'peoplegroups.org', 'unhcr.org', '28toomany.org', 'pewforum.org', 'unhcr.org', 'unhcr.org', 'www.mises.org', ['plos genetics'], ['nature'], [' american journal of human genetics '], ['molecular biology and evolution'], ['scientific reports '], ['springer'], [' bmc genomics '], ['the american journal of human genetics'], ['european journal of human genetics '], ['scientific reports'], ['annales d'], ['forensic science international'], ['american journal of physical anthropology'], ['annals of human genetics '], ['computers and translation'], ['european journal of human genetics']]",1571696,Require autoconfirmed or confirmed access (no expiry set),153325,5 March 2005,Eleassar777 ,6878,0,2005-03-05,2005-03,2005
345,345,Sri Lankan Tamils,https://en.wikipedia.org/wiki/Sri_Lankan_Tamils,192,11,"['10.2307/2058433', None, '10.1007/bf00157142', '10.1007/bf00963656', '10.1002/ajpa.1330450112', '10.1525/as.1985.25.9.01p0303g', '10.1080/09557570701828592', '10.1080/09584939408719724', '10.1353/anl.2010.0021', '10.2307/2058432', None, '8543296', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None]","[['[[the journal of asian studies'], ['human biology '], ['[[indo-iranian journal'], ['[[indo-iranian journal'], ['american journal of physical anthropology'], ['[[asian survey'], ['[[cambridge review of international affairs'], ['contemporary south asia'], ['anthropological linguistics'], ['[[journal of asian studies']]",18,9,0,55,0,6,93,0.09375,0.046875,0.2864583333333333,0.057291666666666664,0.0,0.19791666666666666,10,"['www.state.gov', 'www.nas.gov', 'lcweb2.loc.gov', 'www.statistics.gov', 'www.statistics.gov', 'www.statistics.gov', 'www.statistics.gov', 'statistics.gov', 'www.slelections.gov', 'www.tamilnet.com', 'books.google.com', 'www.krepublishers.com', 'books.google.com', 'www.thestar.com', 'www.colombotelegraph.com', 'books.google.com', 'books.google.com', 'books.google.com', 'socialaffairsjournal.com', 'books.google.com', 'frontline.thehindu.com', 'books.google.com', 'economictimes.indiatimes.com', 'books.google.com', 'books.google.com', 'www.newindianexpress.com', 'www.boston.com', 'gateway.proquest.com', 'salem-news.com', 'www.hindu.com', 'tamilculture.com', 'www.colombotelegraph.com', 'books.google.com', 'www.time.com', 'www.hindu.com', 'books.google.com', 'books.google.com', 'www.hindu.com', 'books.google.com', 'www.torontosun.com', 'books.google.com', 'www.ft.com', 'books.google.com', 'frontline.thehindu.com', 'www.theglobeandmail.com', 'books.google.com', 'www.forbes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'glbtq.com', 'www.ejvs.laurasianacademy.com', 'www.google.com', 'www.nationmultimedia.com', 'www.thestar.com', 'www.google.com', 'books.google.com', 'www.bbc.com', 'www.tamilnet.com', 'www.hindu.com', 'articles.timesofindia.indiatimes.com', 'books.google.com', 'www.defonseka.com', 'mahavamsa.org', 'www.jstor.org', 'www.amnesty.org', 'www.eff.org', 'vedda.org', 'www.un.org', 'tamilelibrary.org', 'www.crisisgroup.org', 'murugan.org', 'www.amnesty.org', 'www.satp.org', 'report2007.amnesty.org', 'www.crisisgroup.org', 'archive.ifla.org', 'www.pluralism.org', 'pewforum.org', 'www.ifla.org', 'www.amnesty.org', ['[[the journal of asian studies'], ['human biology '], ['[[indo-iranian journal'], ['[[indo-iranian journal'], ['american journal of physical anthropology'], ['[[asian survey'], ['[[cambridge review of international affairs'], ['contemporary south asia'], ['anthropological linguistics'], ['[[journal of asian studies']]",4096004,Allow all users (no expiry set),123734,16 February 2006,Kanatonian ,3880,26,2006-02-16,2006-02,2006
346,346,Culture of Iran,https://en.wikipedia.org/wiki/Culture_of_Iran,93,8,"['10.1006/jasc.1999.0555', '10.2307/350454', '10.1073/pnas.111163198', '10.1038/444022a', '10.1073/pnas.0801317105', '10.1126/science.290.5496.1485', '10.22059/jfadram.2012.24776', '10.1126/science.287.5461.2254', None, None, '11344280', '17080057', '18697943', '17771221', None, '10731145', None, None, '33220', None, '2575338', None, None, None]","[['  journal of archaeological science'], ['journal of marriage and family'], ['  proceedings of the national academy of sciences'], ['nature'], ['  proceedings of the national academy of sciences'], ['science', 'sciencemag.org'], ['honarhay-e ziba'], [' science ']]",10,1,0,20,0,0,54,0.10752688172043011,0.010752688172043012,0.21505376344086022,0.08602150537634409,0.0,0.20430107526881722,8,"['cia.gov', 'www.nasehpour.com', 'www.krysstal.com', 'www.dw.com', 'about.com', 'ethnologue.com', 'www.ethnologue.com', 'artira.com', 'www.nationmaster.com', 'farsinet.com', 'www.laurelvictoriagray.com', 'www.iran-daily.com', 'www.sairamtour.com', 'www.free-definition.com', 'www.csmonitor.com', 'thebestofhabibi.com', 'www.nytimes.com', 'www.birdnature.com', 'farsinet.com', 'www.forbes.com', 'www.britannica.com', 'whc.unesco.org', 'www.iranicaonline.org', 'www.iranicaonline.org', 'www.iranicaonline.org', 'ungei.org', 'www.iranicaonline.org', 'livius.org', 'www.iran-heritage.org', 'libmma.contentdm.oclc.org', 'www.iranicaonline.org', ['  journal of archaeological science'], ['journal of marriage and family'], ['  proceedings of the national academy of sciences'], ['nature'], ['  proceedings of the national academy of sciences'], ['science', 'sciencemag.org'], ['honarhay-e ziba'], [' science ']]",965233,Allow all users (no expiry set),66539,7 September 2004,Mnamiri ,1496,7,2004-09-07,2004-09,2004
347,347,Nantes,https://en.wikipedia.org/wiki/Nantes,184,4,"['10.1002/joc.3552', '10.1127/0941-2948/2010/0430', '10.1080/00221344508986498', '10.4000/cybergeo.23155', None, None, None, None, None, None, None, None]","[['international journal of climatology '], ['meteorologische zeitschrift '], ['[[journal of geography'], ['cybergeo ']]",5,6,0,31,0,0,139,0.02717391304347826,0.03260869565217391,0.16847826086956522,0.021739130434782608,0.0,0.08152173913043478,4,"['ftp.atdd.noaa.gov', 'seattle.gov', 'www.durban.gov', 'ftp.atdd.noaa.gov', 'www.tbilisi.gov', 'www.cardiff.gov', 'www.nantes-tourisme.com', 'www.collinsdictionary.com', 'www.completefrance.com', 'www.linternaute.com', 'books.google.com', 'www.bbc.com', 'www.nantes-usa.com', 'cdn.ter.sncf.com', 'www.moovitapp.com', 'club-presse-nantes.com', 'www.nantes-developpement.com', 'www.moovitapp.com', 'www.britannica.com', 'www.meteofrance.com', 'www.economist.com', 'club-presse-nantes.com', 'books.google.com', 'www.royal-de-luxe.com', 'medias.sncf.com', 'www.nantes-developpement.com', 'en.oxforddictionaries.com', 'books.google.com', 'nantes.maville.com', 'www.airbusgroup.com', 'rankings.ft.com', 'www.meteofrance.com', 'books.google.com', 'club-presse-nantes.com', 'books.google.com', 'www.telenantes.com', 'www.euronantes.com', 'kr.ambafrance.org', 'creativecommons.org', 'www.loire-estuaire.org', 'www.amtuir.org', 'www.loire-estuaire.org', ['international journal of climatology '], ['meteorologische zeitschrift '], ['[[journal of geography'], ['cybergeo ']]",67453,Allow all users (no expiry set),159008,4 August 2002,Erwan~enwiki ,2442,1,2002-08-04,2002-08,2002
348,348,Luffa,https://en.wikipedia.org/wiki/Luffa,15,6,"['10.1038/162576b0', '10.1016/j.jbiomech.2014.02.010', '10.1016/j.jbiomech.2004.09.027', '10.1016/j.ijimpeng.2013.01.004', '10.1016/j.jmbbm.2012.07.004', None, None, None, None, None, None, None, None, None, None]","[['nature '], ['journal of biomechanics'], ['journal of biomechanics'], ['international journal of impact engineering'], ['journal of the mechanical behavior of biomedical materials']]",0,0,0,7,0,0,2,0.0,0.0,0.4666666666666667,0.4,0.0,0.4,5,"['www.rolexawards.com', 'floridata.com', 'books.google.com', 'www.rumicooks.com', 'www.rumicooks.com', 'udupi-recipes.com', 'www.saffrontrail.com', ['nature '], ['journal of biomechanics'], ['journal of biomechanics'], ['international journal of impact engineering'], ['journal of the mechanical behavior of biomedical materials']]",80993,Allow all users (no expiry set),21471,5 September 2002,PierreAbbat ,739,0,2002-09-05,2002-09,2002
349,349,Thessaloniki,https://en.wikipedia.org/wiki/Thessaloniki,323,1,"['10.1017/s001781600002530x', None, None]",[['harvard theological review']],15,3,0,108,0,0,197,0.04643962848297214,0.009287925696594427,0.33436532507739936,0.0030959752321981426,0.0,0.058823529411764705,1,"['www.ngdc.noaa.gov', 'government.gov', 'earthquake.usgs.gov', 'books.google.com', 'topuniversities.com', 'www.lonelyplanet.com', 'lonelyplanet.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.ekathimerini.com', 'www.eventsinteractive.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thenationalherald.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.greece-is.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.myjewishlearning.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.wewantapplegreece.com', 'books.google.com', 'books.google.com', 'www.tnr.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.yougoculture.com', 'books.google.com', 'books.google.com', 'books.google.com', 'hotelrotonda.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'galanissportsdata.com', 'books.google.com', 'books.google.com', 'travel.nationalgeographic.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.weatherbase.com', 'books.google.com', 'www.greekstatemuseum.com', 'books.google.com', 'books.google.com', 'visitthessalonikigreece.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.ypodomes.com', 'www.worldclimate.com', 'books.google.com', 'books.google.com', 'leicaliker.com', 'issuu.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.haaretz.com', 'books.google.com', 'www.nikiforidis-cuomo.com', 'www.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'galanissportsdata.com', 'www.ypodomes.com', 'books.google.com', 'homelessmontresor.blogspot.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thessalonikibookfair.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.memorialmuseums.org', 'www.worldhistory.org', 'whc.unesco.org', 'www.lpth.org', 'www.olympic.org', 'www.ushmm.org', 'www.promacedonia.org', 'encyclopedia.ushmm.org', 'www.alexanderthegreatmarathon.org', 'mmca.org', 'en.climate-data.org', 'www.worldclimate.org', 'wikimapia.org', 'www.seegames2007.org', 'www.lpth.org', ['harvard theological review']]",40471,Allow all users (no expiry set),250852,19 October 2001,216.99.203.xxx ,7469,3,2001-10-19,2001-10,2001
350,350,Pontic Greeks,https://en.wikipedia.org/wiki/Pontic_Greeks,147,8,"['10.2307/631221', '10.2307/3642433', 'abs/10.4133/1.4721889', '10.2307/1845120', '10.4305/metu.jfa.2012.1.14', '10.4000/anatoli.315', '10.2307/1291371', None, None, None, None, None, None, None, None, None, None, None, None, None, None]","[[' the journal of hellenic studies'], ['anatolian studies '], ['symposium on the application of geophysics to engineering and environmental problems 2012 '], ['the american historical review ', 'oxford university press'], ['metu journal of the faculty of architecture '], ['[[anatoli '], ['dumbarton oaks papers ']]",9,11,0,54,0,0,65,0.061224489795918366,0.07482993197278912,0.3673469387755102,0.05442176870748299,0.0,0.19047619047619047,7,"['www.sinop.adalet.gov', 'www.rizekulturturizm.gov', 'giresun.ktb.gov', 'gumushane.gov', 'www.sebinkarahisar.gov', 'www.kulturportali.gov', 'www.sumela.gov', 'kvmgm.ktb.gov', 'www.giresun.gov', 'sinop.ktb.gov', 'giresun.ktb.gov', 'www.google.com', 'books.google.com', 'imdb.com', 'pontosworld.com', 'www.google.com', 'pontosworld.com', 'books.google.com', 'angelfire.com', 'www.youtube.com', 'www.google.com', 'imdb.com', 'karalahana.com', 'books.google.com', 'www.karalahana.com', 'karalahana.com', 'pontosworld.com', 'www.dailysabah.com', 'www.youtube.com', 'tr.blackseasilkroad.com', 'www.google.com', 'pontosworld.com', 'imdb.com', 'www.karalahana.com', 'www.bbc.com', 'www.haberler.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.google.com', 'www.hurriyetdailynews.com', 'books.google.com', 'www.dimiourgiestisnias.com', 'books.google.com', 'www.aa.com', 'imdb.com', 'www.karalahana.com', 'pontosworld.com', 'imdb.com', 'peristereota.com', 'www.google.com', 'imdb.com', 'www.google.com', 'www.britannica.com', 'www.ijhssnet.com', 'imturkey.com', 'pontosworld.com', 'www.google.com', 'www.huffpost.com', 'pontosworld.com', 'www.google.com', 'www.karalahana.com', 'pontosworld.com', 'journals.openedition.org', 'turkiyekulturvarliklari.hrantdink.org', 'www.jstor.org', 'www.jstor.org', 'www.worldhistory.org', 'dergipark.org', 'whc.unesco.org', 'en.wikisource.org', 'whc.unesco.org', [' the journal of hellenic studies'], ['anatolian studies '], ['symposium on the application of geophysics to engineering and environmental problems 2012 '], ['the american historical review ', 'oxford university press'], ['metu journal of the faculty of architecture '], ['[[anatoli '], ['dumbarton oaks papers ']]",1619567,Allow all users (no expiry set),98123,18 March 2005,Briangotts ,1504,14,2005-03-18,2005-03,2005
351,351,Kolhapur,https://en.wikipedia.org/wiki/Kolhapur,42,0,[],[],0,6,0,32,0,0,4,0.0,0.14285714285714285,0.7619047619047619,0.0,0.0,0.14285714285714285,0,"['mahasdb.maharashtra.gov', 'www.kolhapurcorporation.gov', 'imdpune.gov', 'cultural.maharashtra.gov', 'imdpune.gov', 'www.kolhapurcorporation.gov', 'books.google.com', 'books.google.com', 'maharashtratimes.indiatimes.com', 'archive.indianexpress.com', 'www.thehindu.com', 'books.google.com', 'maharashtratimes.indiatimes.com', 'prabhupadabooks.com', 'archive.indianexpress.com', 'books.google.com', 'www.reportagebygettyimages.com', 'books.google.com', 'm.maharashtratimes.com', 'www.ambabai.com', 'books.google.com', 'books.google.com', 'maharashtratimes.indiatimes.com', 'ibnlive.in.com', 'maps.google.com', 'books.google.com', 'maharashtratimes.indiatimes.com', 'www.business-standard.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'economictimes.indiatimes.com', 'www.demographia.com', 'timesofindia.indiatimes.com', 'www.sacred-texts.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'land.com']",337536,Allow all users (no expiry set),40932,9 October 2003,Maheshkale ,3732,14,2003-10-09,2003-10,2003
352,352,Malabar District,https://en.wikipedia.org/wiki/Malabar_District,112,2,"['10.2307/2690896', '10.1086/356288', None, None, None, None]","[['mathematics magazine '], ['isis ']]",4,17,0,34,0,0,55,0.03571428571428571,0.15178571428571427,0.30357142857142855,0.017857142857142856,0.0,0.20535714285714285,2,"['lsi.gov', 'lsi.gov', 'lsi.gov', 'lsi.gov', 'dmg.kerala.gov', 'lsi.gov', 'lsi.gov', 'lsi.gov', 'lsi.gov', 'censusindia.gov', 'censusindia.gov', 'legislative.gov', 'mahe.gov', 'lsi.gov', 'lsi.gov', 'censusindia.gov', 'lsi.gov', 'ananthapuri.com', 'books.google.com', 'books.google.com', 'www.facesplacesandplates.com', 'books.google.com', 'books.google.com', 'www.deccanchronicle.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'www.thehindu.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.asianage.com', 'www.thehindu.com', 'www.cookawesome.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'www.thetakeiteasychef.com', 'frontline.thehindu.com', 'books.google.com', 'dcbookstore.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.hindu.com', 'books.google.com', 'books.google.com', 'www.cartage.org', 'www.gutenberg.org', 'www.worldstatesmen.org', 'www.cpimkerala.org', ['mathematics magazine '], ['isis ']]",3563411,Require administrator access (no expiry set),150757,29 December 2005,Tom Radulovich ,717,0,2005-12-29,2005-12,2005
353,353,North Rhine-Westphalia,https://en.wikipedia.org/wiki/North_Rhine-Westphalia,37,0,[],[],4,0,0,5,0,0,28,0.10810810810810811,0.0,0.13513513513513514,0.0,0.0,0.10810810810810811,0,"['www.kitchenproject.com', 'de.statista.com', 'www.neweuropeaneconomy.com', 'www.oeffnungszeiten.com', 'de.statista.com', 'en.wikipedia.org', 'hdi.globaldatalab.org', 'hdi.globaldatalab.org', 'www.eurofir.org']",38414,Allow all users (no expiry set),70445,17 May 2001,LA2 ,1581,7,2001-05-17,2001-05,2001
354,354,Saxony,https://en.wikipedia.org/wiki/Saxony,35,0,[],[],2,0,0,5,0,0,28,0.05714285714285714,0.0,0.14285714285714285,0.0,0.0,0.05714285714285714,0,"['www.economist.com', 'gurdwara-germany.com', 'www.washingtonpost.com', 'www.deseretnews.com', 'de.statista.com', 'hdi.globaldatalab.org', 'www.churchofengland.org']",28395,Allow all users (no expiry set),66986,17 May 2001,LA2 ,1466,5,2001-05-17,2001-05,2001
355,355,Qing dynasty,https://en.wikipedia.org/wiki/Qing_dynasty,138,18,"['10.1215/01636545-2004-88-193', '10.2307/2659026', '10.1177/0097700405282349', '10.2307/2646525', '10.1080/1547402x.2016.1168180', '10.2307/2051924', '10.1111/0020-8833.00053', '10.1017/s0021911800022713', '10.2307/2645062', '10.1111/j.1467-8306.1979.tb01285.x', '10.1111/j.1478-0542.2012.00841.x', '10.2753/csh0009-4633430208', '10.2307/2718931', '10.2307/2658945', '10.1891/1062-8061.4.1.129', '10.1111/j.1754-0208.2011.00454.x', '10.1017/s0026749x00005333', '10.2307/2056359', None, None, None, None, None, None, None, None, None, None, None, None, None, None, '7581277', None, None, '11617269', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None]","[[' radical history review '], [' the journal of asian studies '], [' modern china '], [' the journal of asian studies '], ['chinese historical review'], [' the journal of asian studies '], ['[[international studies quarterly'], ['journal of asian studies'], ['asian survey'], ['annals of the association of american geographers'], ['history compass'], ['chinese studies in history '], [' harvard journal of asiatic studies '], [' [[journal of asian studies'], ['nursing history review'], [' journal for eighteenth-century studies '], ['modern asian studies'], ['journal of asian studies']]",4,0,0,37,0,0,79,0.028985507246376812,0.0,0.26811594202898553,0.13043478260869565,0.0,0.15942028985507245,18,"['books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'gotheborg.com', 'books.google.com', 'books.google.com', 'brill.com', 'www.berkshirepublishing.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'wayoftheeating.wordpress.com', 'www.lingnanart.com', 'www.scmp.com', 'www.britannica.com', 'www.google.com', 'books.google.com', 'timesmachine.nytimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.google.com', 'books.google.com', 'china.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'www.artsmia.org', 'www.danwei.org', 'www.metmuseum.org', 'escholarship.org', [' radical history review '], [' the journal of asian studies '], [' modern china '], [' the journal of asian studies '], ['chinese historical review'], [' the journal of asian studies '], ['[[international studies quarterly'], ['journal of asian studies'], ['asian survey'], ['annals of the association of american geographers'], ['history compass'], ['chinese studies in history '], [' harvard journal of asiatic studies '], [' [[journal of asian studies'], ['nursing history review'], [' journal for eighteenth-century studies '], ['modern asian studies'], ['journal of asian studies']]",25310,Require administrator access (no expiry set),168694,20 November 2001,Chenyu ,7993,19,2001-11-20,2001-11,2001
356,356,Kannur district,https://en.wikipedia.org/wiki/Kannur_district,60,0,[],[],5,15,0,22,0,0,18,0.08333333333333333,0.25,0.36666666666666664,0.0,0.0,0.3333333333333333,0,"['censusindia.gov', 'kannur.keralapolice.gov', 'mahe.gov', 'censusindia.gov', 'www.ecostat.kerala.gov', 'www.censusindia.gov', 'censusindia.gov', 'www.censusindia.gov', 'ceo.kerala.gov', 'censusindia.gov', 'www.dic.kerala.gov', 'sec.kerala.gov', 'www.censusindia.gov', 'lsi.gov', 'censusindia.gov', 'books.google.com', 'www.thehindu.com', 'www.deccanchronicle.com', 'ananthapuri.com', 'www.thehindu.com', 'www.arabnews.com', 'www.deccanherald.com', 'www.thetakeiteasychef.com', 'books.google.com', 'www.thenewsminute.com', 'books.google.com', 'books.google.com', 'www.deccanchronicle.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.thehindu.com', 'www.facesplacesandplates.com', 'www.bbc.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.keralaculture.org', 'www.kottayamad.org', 'keralafolklore.org', 'www.keralatourism.org', 'www.in.undp.org']",865032,Require administrator access (no expiry set),53912,29 July 2004,Sreejith p menon ,1816,7,2004-07-29,2004-07,2004
357,357,Tibet,https://en.wikipedia.org/wiki/Tibet,133,6,"['10.16249/j.cnki.1005-5738.2007.02.006', '10.1007/s12231-008-9038-3', '10.1146/annurev-animal-021815-111155', '10.1073/pnas.0907844106', None, None, '26526544', '19955425', None, None, None, '2795552']","[['journal of tibet university '], ['economic botany'], ['[[annual review of animal biosciences', '[[annual reviews '], [' proc natl acad sci u s a ']]",11,11,0,26,0,1,79,0.08270676691729323,0.08270676691729323,0.19548872180451127,0.045112781954887216,0.0,0.21052631578947367,4,"['www.cia.gov', 'old-cdc.cma.gov', 'www.neac.gov', 'www.imd.gov', 'www.xzta.gov', 'www.cia.gov', 'oceanservice.noaa.gov', 'www.eng.yn.gov', 'www.mausam.gov', 'webarchive.loc.gov', 'www.uscirf.gov', 'english.people.com', 'www.religionfacts.com', 'ogimet.com', 'www.france24.com', 'news.xinhuanet.com', 'articles.latimes.com', 'books.google.com', 'www.bbc.com', 'www.nytimes.com', 'science.nationalgeographic.com', 'books.google.com', 'books.google.com', 'www.tibet.com', 'books.google.com', 'books.google.com', 'sites.google.com', 'books.google.com', 'query.nytimes.com', 'news.xinhuanet.com', 'thediplomat.com', 'voyage.typepad.com', 'books.google.com', 'bloomberg.com', 'www.nytimes.com', 'sites.google.com', 'www.tibetlink.com', 'www.refworld.org', 'www.npr.org', 'tew.org', 'stason.org', 'www.globalsecurity.org', 'www.mherrera.org', 'www.eastwestcenter.org', 'www.eastwestcenter.org', 'www.eastwestcenter.org', 'circleofblue.org', 'www.tibetjustice.org', ['journal of tibet university '], ['economic botany'], ['[[annual review of animal biosciences', '[[annual reviews '], [' proc natl acad sci u s a ']]",31516,Require administrator access (no expiry set),110729,12 January 2002,152.163.197.xxx ,8166,11,2002-01-12,2002-01,2002
358,358,Syria,https://en.wikipedia.org/wiki/Syria,275,9,"['10.1080/07075332.2017.1367705', '10.1038/s41467-020-19493-3', '10.1093/biosci/bix014', '10.1080/00263208908700793', '10.1086/511103', '10.1086/373570', '10.1086/374384', None, '33293507', '28608869', None, None, None, '12629598', None, '7723057', '5451287', None, None, None, '1180338']","[['the international history review'], ['nature communications'], ['bioscience'], ['middle eastern studies'], [' journal of near eastern studies '], [' journal of near eastern studies '], ['american journal of human genetics ']]",42,12,0,125,0,7,80,0.15272727272727274,0.04363636363636364,0.45454545454545453,0.03272727272727273,0.0,0.2290909090909091,7,"['state.gov', 'state.gov', '2009-2017.state.gov', 'www.mohe.gov', 'ste.gov', '2009-2017.state.gov', 'www.mohe.gov', 'www.cia.gov', 'hwb.gov', 'mofa.gov', 'www.cia.gov', 'moct.gov', 'www.scribd.com', 'books.google.com', 'uk.reuters.com', 'books.google.com', 'www.haaretz.com', 'www.jpost.com', 'www.nytimes.com', 'www.nytimes.com', 'www.time.com', 'www.nytimes.com', 'edition.cnn.com', 'books.google.com', 'www.nytimes.com', 'www.fw-magazine.com', 'global.oup.com', 'www.newspapers.com', 'news.yahoo.com', 'www.reuters.com', 'www.wsj.com', 'www.aljazeera.com', 'www.al-monitor.com', 'everything2.com', 'www.torontosun.com', 'euronews.com', 'www.washingtonpost.com', 'www.etymonline.com', 'news.yahoo.com', 'www.dailystar.com', 'books.google.com', 'naharnet.com', 'www.fw-magazine.com', 'www.nytimes.com', 'www.jpost.com', 'www.huffingtonpost.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.newsweek.com', 'books.google.com', 'www.dailystar.com', 'www.worldatlas.com', 'www.ynetnews.com', 'ancienthistory.about.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'www.reuters.com', 'ancientneareast.tripod.com', 'www.scribd.com', 'www.todayszaman.com', 'www.fw-magazine.com', 'books.google.com', 'news24.com', 'www.ft.com', 'www.bbc.com', 'www.newspapers.com', 'www.britannica.com', 'books.google.com', 'www.foxnews.com', 'magma.nationalgeographic.com', 'www.cnn.com', 'www.reuters.com', 'www.nytimes.com', 'www.arabnews.com', 'www.syriauntold.com', 'books.google.com', 'books.google.com', '2fwww.theglobeandmail.com', 'books.google.com', 'books.google.com', 'www.theglobeandmail.com', 'books.google.com', 'www.scribd.com', 'www.chinadaily.com', 'www.reuters.com', 'www.scribd.com', 'www.reuters.com', 'books.google.com', 'www.usatoday.com', 'edition.cnn.com', 'books.google.com', 'books.google.com', 'www.israelnationalnews.com', 'www.reuters.com', 'www.slate.com', 'forward.com', 'books.google.com', 'www.fw-magazine.com', 'books.google.com', 'www.google.com', 'www.arabnews.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'www.ft.com', 'www.indexmundi.com', 'books.google.com', 'www.usatoday.com', 'www.algemeiner.com', 'www.syriahr.com', 'books.google.com', 'books.google.com', 'www.france24.com', '2fwww.theglobeandmail.com', 'www.saudiaramcoworld.com', 'www.newsweek.com', 'www.britannica.com', 'www.cnn.com', 'www.scribd.com', 'www.nytimes.com', 'www.nytimes.com', 'www.foreignaffairs.com', 'news.xinhuanet.com', 'books.google.com', 'www.ft.com', 'www.vice.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'www.etymonline.com', 'books.google.com', 'books.google.com', 'www.goshennews.com', 'seat61.com', 'www.jewishvirtuallibrary.org', 'www.hrw.org', 'www.carnegieendowment.org', 'www.jaas.org', 'carnegieendowment.org', 'www.freedomhouse.org', 'www.ohchr.org', 'www.data.unhcr.org', 'www.sesrtcic.org', 'www.hrw.org', 'www.jaas.org', 'www-wds.worldbank.org', 'freedomhouse.org', 'data.worldbank.org', 'globalsecurity.org', 'visionofhumanity.org', 'www.refugees.org', 'www.metmuseum.org', 'hosted2.ap.org', 'metmuseum.org', 'freedomhouse.org', 'siteresources.worldbank.org', 'www.data.unhcr.org', 'www.unhcr.org', 'documents1.worldbank.org', 'www.unhcr.org', 'www.unhcr.org', 'hdr.undp.org', 'www.witness-pioneer.org', 'data.worldbank.org', 'ftp.fao.org', 'population.un.org', 'www.carnegieendowment.org', 'siteresources.worldbank.org', 'www.ilo.org', 'www.data.unhcr.org', 'www.fearab.org', 'www.heritage.org', 'www.meforum.org', 'www.impact-se.org', 'www.sesrtcic.org', 'golan-marsad.org', ['the international history review'], ['nature communications'], ['bioscience'], ['middle eastern studies'], [' journal of near eastern studies '], [' journal of near eastern studies '], ['american journal of human genetics ']]",7515849,Require administrator access (no expiry set),184990,28 May 2001,KoyaanisQatsi ,10044,26,2001-05-28,2001-05,2001
359,359,Catalonia,https://en.wikipedia.org/wiki/Catalonia,213,5,"['10.1016/j.jhevol.2005.10.001', '10.2307/337523', '10.1111/imig.12323', '10.3406/ecelt.1948.1196', '16364406', None, None, None, None, None, None, None]","[[' journal of human evolution '], ['hispania '], ['international migration'], ['études celtiques']]",9,2,0,64,0,3,130,0.04225352112676056,0.009389671361502348,0.3004694835680751,0.023474178403755867,0.0,0.07511737089201878,4,"['soir.senate.ca.gov', 'soir.senate.ca.gov', 'noticias.juridicas.com', 'www.economist.com', 'www.thetrainline.com', 'lavanguardia.com', 'www.elpais.com', 'books.google.com', 'ethnologue.com', 'es.opinometre.com', 'noticias.juridicas.com', 'cadenaser.com', 'books.google.com', 'www.lavanguardia.com', 'www.britannica.com', 'blogs.periodistadigital.com', 'costabravatouristguide.com', 'books.google.com', 'www.lavanguardia.com', 'www.bbc.com', 'books.google.com', 'publimetro.com', 'www.info7.com', 'world.time.com', 'books.google.com', 'www.antena3.com', 'datosmacro.com', 'www.elperiodico.com', 'books.google.com', 'www.bergueda.com', 'www.thetrainline.com', 'www.datosmacro.com', 'www.demographia.com', 'economist.com', 'news.scotsman.com', 'www.washingtonpost.com', 'www.cnbc.com', 'www.reuters.com', 'elpais.com', 'books.google.com', 'elpais.com', 'euobserver.com', 'www.lavanguardia.com', 'noticias.juridicas.com', 'blogs.periodistadigital.com', 'etymonline.com', 'articles.economictimes.indiatimes.com', 'www.lavanguardia.com', 'elpais.com', 'books.google.com', 'cava-and-co.com', 'www.expatica.com', 'www.fira-aer-rugby.com', 'racalacarta.com', 'www.expansion.com', 'books.google.com', 'www.youtube.com', 'books.google.com', 'www.libremercado.com', 'www.railwaygazette.com', 'www.railjournal.com', 'books.google.com', 'expansión.com', 'www.elpais.com', 'www.bloomberg.com', 'books.google.com', 'wayback.archive-it.org', 'www.histoire-empire.org', 'www.pbs.org', 'hdi.globaldatalab.org', 'unpo.org', 'www.edmaktub.org', 'www.imf.org', 'www.histoire-empire.org', 'europeanregionofgastronomy.org', [' journal of human evolution '], ['hispania '], ['international migration'], ['études celtiques']]",6822,Allow all users (no expiry set),198829,17 October 2001,Tsja ,8006,17,2001-10-17,2001-10,2001
360,360,Chios,https://en.wikipedia.org/wiki/Chios,54,2,"['10.5194/nhess-5-717-2005', None, None]",[['natural hazards and earth system sciences ']],6,0,0,5,0,0,41,0.1111111111111111,0.0,0.09259259259259259,0.037037037037037035,0.0,0.14814814814814814,1,"['www.com', 'dictionary.com', 'books.google.com', 'www.firstworldwar.com', 'www.ancientlibrary.com', 'www.livius.org', 'chianfed.org', 'sephardicstudies.org', 'livius.org', 'www.greece.org', 'www.eoearth.org', ['natural hazards and earth system sciences ']]",17067,Allow all users (no expiry set),49268,25 February 2002,Conversion script ,1597,6,2002-02-25,2002-02,2002
361,361,Tirupati,https://en.wikipedia.org/wiki/Tirupati,116,0,[],[],14,20,0,67,0,0,15,0.1206896551724138,0.1724137931034483,0.5775862068965517,0.0,0.0,0.29310344827586204,0,"['www.aptdc.gov', 'www.portal.gsi.gov', 'cdma.gov', 'imdpune.gov', 'www.appolice.gov', 'imdpune.gov', 'city.imd.gov', 'www.indianrailways.gov', 'mct.gov', 'census.gov', 'censusindia.gov', 'censusindia.gov', 'tirupati.cdma.ap.gov', 'www.censusindia.gov', 'www.tuda.gov', 'www.tuda.gov', 'www.aptdc.gov', 'aproads.cgg.gov', 'www.ap.gov', 'www.portal.gsi.gov', 'www.thehindu.com', 'daily.bhaskar.com', 'www.deccanchronicle.com', 'www.thehindu.com', 'www.newindianexpress.com', 'www.business-standard.com', 'books.google.com', 'www.thehindu.com', 'www.deccanherald.com', 'economictimes.indiatimes.com', 'books.google.com', 'www.thehindubusinessline.com', 'www.youtube.com', 'www.thehindu.com', 'indianexpress.com', 'www.newindianexpress.com', 'indianexpress.com', 'www.thehindu.com', 'books.google.com', 'www.thehindu.com', 'www.newindianexpress.com', 'www.geocities.com', 'www.newindianexpress.com', 'www.thehindubusinessline.com', 'www.india.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehansindia.com', 'www.uniindia.com', 'www.thehansindia.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehindu.com', 'books.google.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehindubusinessline.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.thehindu.com', 'india.com', 'economictimes.indiatimes.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehindubusinessline.com', 'www.youtube.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.thehindu.com', 'books.google.com', 'www.thehansindia.com', 'www.eco-web.com', 'www.newindianexpress.com', 'www.ndtv.com', 'www.siasat.com', 'www.thehindu.com', 'www.newindianexpress.com', 'www.thehindu.com', 'www.thehindu.com', 'www.newindianexpress.com', 'www.tirupaticorporation.org', 'www.tirumala.org', 'www.birrd.org', 'www.tirumala.org', 'www.tirupaticorporation.org', 'www.tirumala.org', 'svzoo.org', 'www.sangeetasudha.org', 'news.tirumala.org', 'ttdgoshala.org', 'www.svvedicuniversity.org', 'www.unece.org', 'www.tirumala.org', 'www.tirumala.org']",2892130,Allow all users (no expiry set),75330,12 October 2005,Vyzasatya ,3606,28,2005-10-12,2005-10,2005
362,362,Tallinn,https://en.wikipedia.org/wiki/Tallinn,115,2,"['10.3176/earth.2010.1.03', '10.5194/hess-11-1633-2007', None, None, None, None]","[['estonian journal of earth sciences'], ['hydrol. earth syst. sci. ']]",6,0,0,32,0,1,74,0.05217391304347826,0.0,0.2782608695652174,0.017391304347826087,0.0,0.06956521739130435,2,"['www.copterline.com', 'books.google.com', 'www.copterline.com', 'www.baltictimes.com', 'books.google.com', 'select.nytimes.com', 'books.google.com', 'balticbusinessnews.com', 'books.google.com', 'estonianworld.com', 'encyclopedia2.thefreedictionary.com', 'www.forbes.com', 'books.google.com', 'portoftallinn.com', 'thefreedictionary.com', 'www.airport-business.com', 'techcrunch.com', 'www.kommersant.com', 'www.cushmanwakefield.com', 'www.wsj.com', 'www.arvato.com', 'www.uswitch.com', 'dictionary.infoplease.com', 'books.google.com', 'books.google.com', 'visitestonia.com', 'www.theage.com', 'www.timeanddate.com', 'www.weather-atlas.com', 'visitestonia.com', 'jobs.skype.com', 'books.google.com', 'whc.unesco.org', 'www.easac.org', 'runeberg.org', 'whc.unesco.org', 'www.nonviolent-conflict.org', 'dbs.bh.org', ['estonian journal of earth sciences'], ['hydrol. earth syst. sci. ']]",31577,Allow all users (no expiry set),105604,20 January 2002,Sjc ,3224,24,2002-01-20,2002-01,2002
363,363,Central Europe,https://en.wikipedia.org/wiki/Central_Europe,168,3,"['10.1038/nature.2012.12020', '10.2307/621131', '10.1093/ehr/cej100', None, None, None, None, None, None]","[['nature news '], [' transactions and papers '], ['the english historical review']]",26,6,0,45,0,0,89,0.15476190476190477,0.03571428571428571,0.26785714285714285,0.017857142857142856,0.0,0.20833333333333334,3,"['www.stat.gov', 'www.cia.gov', 'portoncv.gov', 'www.stat.gov', 'stat.gov', 'pod2.stat.gov', 'www.oup.com', 'www.newstatesman.com', 'literalab.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'www.nytimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'centraleuropethrowdown.com', 'highbeam.com', 'www.ebrd.com', 'books.google.com', 'masticationmonologues.com', 'encarta.msn.com', 'timeanddate.com', 'books.google.com', 'books.google.com', 'books.google.com', 'wps.ablongman.com', 'www.newyorker.com', 'www.tholons.com', 'www.railwaypro.com', 'books.google.com', 'www.foreignaffairs.com', 'www.tv.com', 'www.google.com', 'www.oup.com', 'a-ztours.com', 'angelus.com', 'emersonkent.com', 'www.grin.com', 'www.economist.com', 'books.google.com', 'chronicle.com', 'books.google.com', 'books.google.com', 'thefreedictionary.com', 'www.prosperity.com', 'books.google.com', 'www.economist.com', 'www.latimes.com', 'edition.cnn.com', 'hostmonster.com', 'zacat.gesis.org', 'www.ajcarchives.org', 'www.icpdr.org', 'transparency.org', 'www.unhcr-centraleurope.org', 'historyguide.org', 'unstats.un.org', 'science.jrank.org', 'science.jrank.org', 'www.opensocietyfoundations.org', 'science.jrank.org', 'www.ais.unwater.org', 'unstats.un.org', 'w3.unece.org', 'www.visionofhumanity.org', 'www.oecd.org', 'www.transcend.org', 'www.un.org', 'www.rs.undp.org', 'internationaltransportforum.org', 'www.culturelink.org', 'h-net.org', 'www3.weforum.org', 'www.h-net.org', 'faostat3.fao.org', 'centraleurope.org', ['nature news '], [' transactions and papers '], ['the english historical review']]",5188,Allow all users (no expiry set),106774,10 December 2001,Szopen ,4648,13,2001-12-10,2001-12,2001
364,364,Basel,https://en.wikipedia.org/wiki/Basel,119,0,[],[],5,0,0,16,0,0,98,0.04201680672268908,0.0,0.13445378151260504,0.0,0.0,0.04201680672268908,0,"['www.crossair.com', 'www.swiss.com', 'travel.nytimes.com', 'www.ciba.com', 'mobilityexchange.mercer.com', 'saint-louis.plan-interactif.com', 'archives.newyorker.com', 'www.infolignes.com', 'mobilityexchange.mercer.com', 'www.swiss.com', 'www.lifeinbasel.com', 'www.getlisty.com', 'apps2.ubs.com', 'www.basel.com', 'www.weatherbase.com', 'world.com', 'www.bis.org', 'www.bis.org', 'fondationfernet-branca.org', 'www.swissinfo.org', 'www.schaulager.org']",4911,Allow all users (no expiry set),122516,30 December 2001,62.2.17.xxx ,2402,6,2001-12-30,2001-12,2001
365,365,Veneto,https://en.wikipedia.org/wiki/Veneto,90,0,[],[],5,0,0,17,0,1,67,0.05555555555555555,0.0,0.18888888888888888,0.0,0.0,0.05555555555555555,0,"['www.seattlepi.com', 'www.bbc.com', 'www.nytimes.com', 'data.mongabay.com', 'books.google.com', 'www.bbc.com', 'www.collinsdictionary.com', 'query.nytimes.com', 'www.cnn.com', 'www.washingtonpost.com', 'www.adnkronos.com', 'www.nybooks.com', 'adnkronos.com', 'www.raixevenete.com', 'www.wine-searcher.com', 'www.fineartprintsondemand.com', 'www.cbsnews.com', 'whc.unesco.org', 'whc.unesco.org', 'hdi.globaldatalab.org', 'whc.unesco.org', 'whc.unesco.org']",43780,Allow all users (no expiry set),109162,11 March 2002,151.24.146.109 ,2486,1,2002-03-11,2002-03,2002
366,366,Sussex,https://en.wikipedia.org/wiki/Sussex,202,1,"['10.2307/2597413', None, None]",[['economic history review']],28,15,0,20,0,4,134,0.13861386138613863,0.07425742574257425,0.09900990099009901,0.0049504950495049506,0.0,0.21782178217821782,1,"['www.gov', 'scotlandcensus.gov', 'www.ons.gov', 'www.ons.gov', 'www.gov', 'www.southdowns.gov', 'www.eastsussex.gov', 'www.ons.gov', 'www.westsussex.gov', 'www.ons.gov', 'www.metoffice.gov', 'midsussex.gov', 'www.southdowns.gov', 'webarchive.nationalarchives.gov', 'www.statistics.gov', 'techcrunch.com', 'www.ospreypublishing.com', 'www.debretts.com', 'www.oxforddnb.com', 'sussexflag.wordpress.com', 'sussexflag.wordpress.com', 'history-tourist.com', 'www.economist.com', 'www.cricinfo.com', 'historicalfoods.com', 'www.francisfrith.com', 'britannica.com', 'theenglishappleman.com', 'www.thechampagnecompany.com', 'travel.nationalgeographic.com', 'www.topuniversities.com', 'www.economist.com', 'historicalfoods.com', 'www.nytimes.com', 'www.ukrockfestivals.com', 'www.charleston.org', 'www.sussexgiving.org', 'www.ibiblio.org', 'www.dannyhouse.org', 'econjwatch.org', 'www.nobelprize.org', 'www.naturalengland.org', 'www.pallant.org', 'hastingspride.org', 'www.nobelprize.org', 'www.oldpolicecellsmuseum.org', 'www.pbs.org', 'www.prebendalschool.org', 'www.royalsussex.org', 'pallant.org', 'www.scfl.org', 'www.britishmuseum.org', 'www.visitsussex.org', 'www.westdean.org', 'www.sussexrecordsociety.org', 'www.brightonphil.org', 'www.nobelprize.org', 'www.visitsussex.org', 'steyningmuseum.org', 'kipling.org', 'www.fondation-fyssen.org', 'www.nobelprize.org', 'www.theparisreview.org', ['economic history review']]",49699,Allow all users (no expiry set),114345,19 April 2002,Amillar ,1833,12,2002-04-19,2002-04,2002
367,367,Hyderabadi Muslims,https://en.wikipedia.org/wiki/Hyderabadi_Muslims,88,1,"['10.1080/13602008508715945', None, None]","[['journal of muslim minority affairs ', '[[routledge']]",1,1,0,69,0,0,16,0.011363636363636364,0.011363636363636364,0.7840909090909091,0.011363636363636364,0.0,0.03409090909090909,1,"['www.censusindia.gov', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'telanganatoday.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.india-seminar.com', 'books.google.com', 'www.dawn.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.thefridaytimes.com', 'books.google.com', 'www.deccanchronicle.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.news18.com', 'archive.siasat.com', 'www.news18.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.thenewsminute.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'archive.siasat.com', 'www.thenewsminute.com', 'books.google.com', 'www.newindianexpress.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'news.google.com', 'india.blogs.nytimes.com', 'archive.siasat.com', 'archive.siasat.com', 'time.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'archive.siasat.com', 'books.google.com', 'books.google.com', 'archive.siasat.com', 'articles.timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'zeenews.india.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'books.google.com', 'news.dawn.com', 'shareefmp.wordpress.com', 'articles.timesofindia.indiatimes.com', 'books.google.com', 'www.prlog.org', ['journal of muslim minority affairs ', '[[routledge']]",3082906,Allow all users (no expiry set),50278,5 November 2005,Jungli ,1380,1,2005-11-05,2005-11,2005
368,368,Urfa,https://en.wikipedia.org/wiki/Urfa,24,0,[],[],4,1,0,8,0,0,11,0.16666666666666666,0.041666666666666664,0.3333333333333333,0.0,0.0,0.20833333333333334,0,"['www.mgm.gov', 'www.todayszaman.com', 'www.jewishencyclopedia.com', 'c86.tumblr.com', 'books.google.com', 'www.thetorah.com', 'www.sabah.com', 'www.weatherbase.com', 'www.hurriyetdailynews.com', 'arsiv.setav.org', 'www.centropa.org', 'archive.archaeology.org', 'armenian-genocide.org']",285533,Allow all users (no expiry set),31994,31 July 2003,Adam Bishop ,1218,2,2003-07-31,2003-07,2003
369,369,Kurdish culture,https://en.wikipedia.org/wiki/Kurdish_culture,14,1,"['10.4000/ejts.5000', None, None]",[['european journal of turkish studies. social sciences on contemporary turkey']],4,1,0,5,0,0,3,0.2857142857142857,0.07142857142857142,0.35714285714285715,0.07142857142857142,0.0,0.42857142857142855,1,"['cabinet.gov', 'books.google.com', 'books.google.com', 'books.google.com', 'www.adventuressheart.com', 'www.bbc.com', 'thekurdishproject.org', 'thekurdishproject.org', 'thekurdishproject.org', 'bnk.institutkurde.org', ['european journal of turkish studies. social sciences on contemporary turkey']]",3913469,Allow all users (no expiry set),10511,31 January 2006,Diyako ,435,10,2006-01-31,2006-01,2006
370,370,Szczecin,https://en.wikipedia.org/wiki/Szczecin,159,0,[],[],0,6,0,11,0,0,142,0.0,0.03773584905660377,0.06918238993710692,0.0,0.0,0.03773584905660377,0,"['www.gov', 'www.gov', 'bdl.stat.gov', 'bdl.stat.gov', 'www.nationalarchives.gov', 'prezydent2010.pkw.gov', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.weatherbase.com', 'www.halp.com', 'books.google.com', 'books.google.com', 'www.weather-atlas.com', 'www.collinsdictionary.com']",28456,Allow all users (no expiry set),110433,4 October 2001,207.215.86.xxx ,3287,1,2001-10-04,2001-10,2001
371,371,Hanoi,https://en.wikipedia.org/wiki/Hanoi,130,10,"['10.5194/hess-11-1633-2007', '10.1177/0042098011408934', '10.1007/s10624-008-9062-9', '10.1016/j.ssaho.2019.100001', '10.1177/0956247819858019', '10.1002/hyp.8315', 'moi:', '10.1017/9780511998492.002', '10.1080/03050060120043411', '10.5509/2005784559', None, None, None, None, '32704235', None, None, None, None, None, None, None, None, None, '7340485', None, None, None, None, None]","[['hydrol. earth syst. sci. '], ['urban studies'], ['dialectical anthropology'], ['social sciences '], ['environment and urbanization'], ['hydrological processes '], ['asian survey'], ['cambridge university press'], ['comparative education'], ['pacific affairs']]",5,20,0,37,0,0,59,0.038461538461538464,0.15384615384615385,0.2846153846153846,0.07692307692307693,0.0,0.2692307692307692,10,"['thongkehanoi.gov', 'vukuzenzele.gov', 'minsk.gov', 'nchmf.gov', 'thongkehanoi.gov', 'phnompenh.gov', 'hanoi.gov', 'thongkehanoi.gov', 'hanoi.gov', 'www.gso.gov', 'www.gso.gov', 'www.monre.gov', 'www.hanoi.gov', 'www.gso.gov', 'www.monre.gov', 'statehouse.gov', 'beijing.gov', 'www.gso.gov', 'thongkehanoi.gov', 'hanoi.gov', 'www.smh.com', 'tnhvietnam.xemzi.com', 'www.businessinsider.com', 'www.restaurants-in-hanoi.com', 'www.theage.com', 'vietnamnews.vnagency.com', 'www.nld.com', '20hanoi.com', 'dotchuoinon.com', 'www.frommers.com', 'visaexplorer.com', 'www.cnn.com', 'www.nytimes.com', 'bbc.com', 'www.vietnamtourism.com', 'www.roughguides.com', 'www.cnn.com', 'global.oup.com', 'www.topuniversities.com', 'www.bbc.com', 'vbusinessnews.com', 'www.com', 'www.f1vietnamgp.com', 'antaranews.com', 'www.willchase.com', 'globalpost.com', 'dantri.com', 'www.thanhniennews.com', 'drive.google.com', 'dantri.com', 'www.formula1.com', 'www.ft.com', 'www.huffingtonpost.com', 'hanoimoi.com', 'smarttravelasia.com', 'www.proquest.com', 'travel.nytimes.com', 'en.unesco.org', 'www.fao.org', 'www2.adb.org', 'www.worldcat.org', 'www.roap.unep.org', ['hydrol. earth syst. sci. '], ['urban studies'], ['dialectical anthropology'], ['social sciences '], ['environment and urbanization'], ['hydrological processes '], ['asian survey'], ['cambridge university press'], ['comparative education'], ['pacific affairs']]",56667,Allow all users (no expiry set),132843,13 June 2002,Zoe ,4039,18,2002-06-13,2002-06,2002
372,372,Dominican Republic,https://en.wikipedia.org/wiki/Dominican_Republic,307,8,"['10.1093/biosci/bix014', '10.2307/978436', '10.1017/s0022050700042182', '10.2307/2546161', '10.1038/s41467-020-19493-3', '10.2747/0272-3646.31.5.455', '10.1017/s0165115300022841', '28608869', None, None, None, '33293507', None, None, '5451287', None, None, None, '7723057', None, None]","[['bioscience'], ['the americas '], [' the journal of economic history'], ['international migration review'], ['nature communications'], ['physical geography '], ['itinerario ']]",52,25,0,125,0,0,98,0.16938110749185667,0.08143322475570032,0.40716612377850164,0.026058631921824105,0.0,0.2768729641693811,7,"['fpc.state.gov', 'www.census.gov', 'ustr.gov', 'ustr.gov', 'factfinder.census.gov', 'lcweb2.loc.gov', 'www.dgii.gov', 'www.bancentral.gov', 'www.cia.gov', 'www.cia.gov', 'www.conapofa.gov', '2009-2017.state.gov', 'www.cia.gov', 'www.seescyt.gov', 'history.state.gov', 'www.cne.gov', 'www.cia.gov', 'www.dgii.gov', 'www.dshs.texas.gov', 'www.conapofa.gov', 'www.dol.gov', 'www.cia.gov', 'history.state.gov', 'cdeee.gov', 'www.senate.gov', 'www.xe.com', 'books.google.com', 'www.reuters.com', 'books.google.com', 'www.eldinero.com', 'sololiteratura.com', 'elnuevodiario.com', 'www.7dias.com', 'www.biografiasyvidas.com', 'www.cielonaranja.com', 'www.diariolibre.com', 'www.laromanabayahibenews.com', 'books.google.com', 'edition.cnn.com', 'www.nytimes.com', 'books.google.com', 'www.britannica.com', 'www.nationsencyclopedia.com', 'xe.com', 'books.google.com', 'books.google.com', 'upi.com', 'books.google.com', 'www.ef.com', 'www.biografiasyvidas.com', 'hoy.com', 'eldia.com', 'www2.dominicantoday.com', 'www.huffingtonpost.com', 'books.google.com', 'diariodigitalrd.com', 'm.diariolibre.com', 'www.topix.com', 'books.google.com', 'www.nytimes.com', 'conectate.com', 'www.cercles.com', 'www.britannica.com', 'www.hispaniola.com', 'www.caribbeannetnews.com', 'www.haitianinternet.com', 'www.nytimes.com', 'dominicantoday.com', 'www.nytimes.com', 'www.smithsonianmag.com', 'www.nytimes.com', 'articles.mcall.com', 'books.google.com', 'encyclopedia.com', 'www.dominicantoday.com', 'acento.com', 'www.nationalgeographic.com', 'books.google.com', 'encarta.msn.com', 'www.7dias.com', 'wcax.com', 'investingnews.com', 'listindiario.com', 'www.dominicantoday.com', 'www.nytimes.com', 'www.elhombrecito.com', 'books.google.com', 'www.listindiario.com', 'books.google.com', 'm.diariolibre.com', 'hoy.com', '7dias.com', 'www.bbc.com', 'listin.com', 'www.abreureport.com', 'huffingtonpost.com', 'books.google.com', 'www.elnuevodiario.com', 'xe.com', 'www.scribd.com', 'content.time.com', 'books.google.com', 'elnacional.com', 'books.google.com', 'video.foxnews.com', 'dominicantoday.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'elnacional.com', 'www.moreorless.au.com', 'www.listindiario.com', 'listin.com', 'www.diariolibre.com', 'books.google.com', 'www.thearda.com', 'biblediscovered.com', 'books.google.com', 'books.google.com', 'www.sobreeldiamante.com', 'www.nytimes.com', 'warfarehistorynetwork.com', 'www.thatsdominican.com', 'books.google.com', 'books.google.com', 'www.sdhoc.com', 'www.bvrd.com', 'nationalgeographic.com', 'elnuevodiario.com', 'www.listindiario.com', 'www.listindiario.com', 'www.listindiario.com', 'xe.com', 'www.diariolibre.com', 'www.colonialzone-dr.com', 'books.google.com', 'dominicanaenmiami.com', 'iasorecords.com', 'xe.com', 'books.google.com', 'books.google.com', 'books.google.com', 'lawrieongold.com', 'books.google.com', 'www.diariolibre.com', 'www.reuters.com', 'www.elcaribe.com', 'www.informejudicial.com', 'www.nytimes.com', 'theworld.org', 'www.centrelink.org', 'www.worldbank.org', 'www.idg.org', 'baseballhall.org', 'www.refworld.org', 'fedojudo.org', 'www.learner.org', 'www.refworld.org', 'www.jewishvirtuallibrary.org', 'www.domrep.org', 'www.dominicanconsulate.org', 'www.oas.org', 'pri.org', 'www.ilo.org', 'whc.unesco.org', 'web.amnesty.org', 'www.jewishvirtuallibrary.org', 'fundacionrenedelrisco.org', 'www.minorityrights.org', 'www.unodc.org', 'www.amnestyusa.org', 'www.globalslaveryindex.org', 'www.weforum.org', 'www.refugeesinternational.org', 'esa.un.org', 'treaties.un.org', 'www.coha.org', 'constitute.org', 'data.worldbank.org', 'www.oas.org', 'www.unesco.org', 'data.worldbank.org', 'whc.unesco.org', 'academiadominicanahistoria.org', 'newsroom.churchofjesuschrist.org', 'www.hrw.org', 'www.wordswithoutborders.org', 'www.worldbank.org', 'unesco.org', 'www.kacike.org', 'www.worldbank.org', 'data.worldbank.org', 'catholictradition.org', 'www.un.org', 'hdr.undp.org', 'data.worldbank.org', 'www.kacike.org', 'www.worldbank.org', 'latinamericanscience.org', 'www.imf.org', 'www.adventistdirectory.org', ['bioscience'], ['the americas '], [' the journal of economic history'], ['international migration review'], ['nature communications'], ['physical geography '], ['itinerario ']]",8060,Require autoconfirmed or confirmed access (no expiry set),259421,5 September 2001,Koyaanis Qatsi ,16224,25,2001-09-05,2001-09,2001
373,373,Gaziantep,https://en.wikipedia.org/wiki/Gaziantep,55,1,"['10.7827/turkishstudies.8598', None, None]",[['international periodical for the languages']],5,3,0,18,0,0,28,0.09090909090909091,0.05454545454545454,0.32727272727272727,0.01818181818181818,0.0,0.16363636363636364,1,"['www.mgm.gov', 'gaziantep.gov', 'minsk.gov', 'www.britannica.com', 'www.endeksa.com', 'books.google.com', 'books.google.com', 'www.milliyet.com', 'www.radikal.com', 'books.google.com', 'www.milliyet.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'www.salom.com', 'books.google.com', 'secim.haberler.com', 'www.britannica.com', 'books.google.com', 'theculturetrip.com', 'books.google.com', 'helenmilesmosaics.org', 'dergipark.org', 'dergipark.org', 'www.ipa-uk.org', 'gso.org', ['international periodical for the languages']]",569037,Allow all users (no expiry set),57385,1 April 2004,TOttenville8 ,1749,2,2004-04-01,2004-04,2004
374,374,Nuremberg,https://en.wikipedia.org/wiki/Nuremberg,68,2,"['10.1016/s0926-6437(99)00014-1', '10.1016/0169-2046(92)90017-t', None, None, None, None]","[['journal of income distribution'], ['landscape and urban planning ']]",2,0,0,14,0,0,50,0.029411764705882353,0.0,0.20588235294117646,0.029411764705882353,0.0,0.058823529411764705,2,"['www.weatherbase.com', 'www.com', 'jewishencyclopedia.com', 'global.oup.com', 'www.airbnb.com', 'www.ricksteves.com', 'www.ricksteves.com', 'www.medievalcoinage.com', 'books.google.com', 'www.com', 'www.ricksteves.com', 'www.thebookseller.com', 'deutsche-pop.com', 'tartanplace.com', 'jwa.org', 'meteo-climat-bzh.dyndns.org', ['journal of income distribution'], ['landscape and urban planning ']]",21287,Allow all users (no expiry set),75189,31 October 2001,H.J. ,2160,13,2001-10-31,2001-10,2001
375,375,Dawoodi Bohra,https://en.wikipedia.org/wiki/Dawoodi_Bohra,210,4,"['10.1093/jis/etr005', '10.1515/islam-2016-0008', '10.15740/has/ajhs/10.1/54-59', None, None, None, None, None, None]","[['journal of islamic studies '], ['der islam'], ['asian journal of home science ']]",15,0,0,146,0,1,44,0.07142857142857142,0.0,0.6952380952380952,0.01904761904761905,0.0,0.09047619047619047,3,"['books.google.com', 'thedawoodibohras.com', 'thedawoodibohras.com', 'www.thehindu.com', 'thedawoodibohras.com', 'tribune.com', 'middleeast.thedawoodibohras.com', 'books.google.com', 'gemsofhistory.com', 'www.thehindubusinessline.com', 'globalnewswire.com', 'books.google.com', 'books.google.com', 'www.thedawoodibohras.com', 'www.chicagotribune.com', 'www.thehindu.com', 'nativeplanet.com', 'www.khaleejtimes.com', 'www.rediff.com', 'mycentraljersey.com', 'www.onmanorama.com', 'sbut.com', 'thedawoodibohras.com', 'timesofindia.indiatimes.com', 'economictimes.indiatimes.com', 'www.khaleejtimes.com', 'usa.thedawoodibohras.com', 'udaipurtimes.com', 'mumbaimirror.indiatimes.com', 'gemsofhistory.com', 'gulfnews.com', 'thedawoodibohras.com', 'www.reuters.com', 'economictimes.indiatimes.com', 'articles.timesofindia.indiatimes.com', 'www.dnaindia.com', 'www.thehindu.com', 'www.khaleejtimes.com', 'malumaat.com', 'www.deccanherald.com', 'books.google.com', 'www.detroitnews.com', 'books.google.com', 'timesofindia.indiatimes.com', 'thedawoodibohras.com', 'sbut.com', 'www.newindianexpress.com', 'thedawoodibohras.com', 'www.indiapost.com', 'books.google.com', 'einnews.com', 'www.thehindu.com', 'www.fnbnews.com', 'teleganatoday.com', 'usa.thedawoodibohras.com', 'timesofindia.indiatimes.com', 'themuslim500.com', 'www.google.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'thedawoodibohras.com', 'globalnewswire.com', 'theroute2roots.com', 'mumbaimirror.indiatimes.com', 'nazafat.com', 'www.thedawoodibohras.com', 'www.thenews.com', 'www.hindustantimes.com', 'www.thedawoodibohras.com', 'gulfnews.com', 'www.journeykitchen.com', 'www.huffpost.com', 'books.google.com', 'usa.thedawoodibohras.com', 'www.sbs.com', 'books.google.com', 'books.google.com', 'books.google.com', 'mumbaimirror.indiatimes.com', 'daijiworld.com', 'www.guinnessworldrecords.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thedawoodibohras.com', 'www.britannica.com', 'www.livemint.com', 'www.straitstimes.com', 'thedawoodibohras.com', 'thedawoodibohras.com', 'indianexpress.com', 'jbasr.com', 'businesswireindia.com', 'economictimes.indiatimes.com', 'www.saifeehospital.com', 'www.business-standard.com', 'thedawoodibohras.com', 'dnaindia.com', 'www.thehindu.com', 'books.google.com', 'thedawoodibohras.com', 'books.google.com', 'www.mumbaifoodie.com', 'ealing.cmis.uk.com', 'thedawoodibohras.com', 'www.khaleejtimes.com', 'books.google.com', 'thedawoodibohras.com', 'www.thehindu.com', 'thedawoodibohras.com', 'uk.thedawoodibohras.com', 'www.thehindu.com', 'canada.thedawoodibohras.com', 'gulfnews.com', 'www.sbut.com', 'economictimes.indiatimes.com', 'www.arabnews.com', 'sbut.com', 'books.google.com', 'food.ndtv.com', 'detroitdawoodibohras.com', 'www.southasia.com', 'www.hindustantimes.com', 'thedawoodibohras.com', 'sbut.com', 'www.straitstimes.com', 'thedawoodibohras.com', 'thedawoodibohras.com', 'nazafat.com', 'www.newindianexpress.com', 'books.google.com', 'www.thenews.com', 'www.smh.com', 'books.google.com', 'www.newindianexpress.com', 'timesofindia.indiatimes.com', 'www.business-standard.com', 'usa.thedawoodibohras.com', 'indianexpress.com', 'www.globenewswire.com', 'mid-day.com', 'mid-day.com', 'finance.yahoo.com', 'islamvoice.com', 'www.thehindu.com', 'escholarship.org', 'www.unicef.org', 'kenyamuseumsociety.org', 'pri.org', 'www.bqhc.org', 'taiseerunnikah.org', 'dronah.org', 'www.manushi-india.org', 'diva-portal.org', 'www.theismaili.org', 'library.oapen.org', 'www.wespeakout.org', 'www.npr.org', 'commons.wikimedia.org', 'www.burhanifoundationindia.org', ['journal of islamic studies '], ['der islam'], ['asian journal of home science ']]",973773,Require autoconfirmed or confirmed access (no expiry set),127818,10 September 2004,203.130.2.98 ,3839,1,2004-09-10,2004-09,2004
376,376,Christmas,https://en.wikipedia.org/wiki/Christmas,281,2,"['10.1162/99608f92.6230ce9f', '10.1093/gmo/9781561592630.article.a2227990', None, None, None, None]","[['harvard data science review'], ['[[grove music online', '[[oxford university press']]",23,4,0,102,0,4,146,0.08185053380782918,0.014234875444839857,0.36298932384341637,0.0071174377224199285,0.0,0.10320284697508897,2,"['www.opm.gov', 'usinfo.state.gov', 'webarchive.loc.gov', 'www.direct.gov', 'books.google.com', 'books.google.com', 'foreignpolicy.com', 'www.britannica.com', 'christianchurchofgod.com', 'citybeat.com', 'www.sacred-destinations.com', 'www.scribd.com', 'www.britannica.com', 'www.bbc.com', 'timetravel-britain.com', 'www.nytimes.com', 'touchstonemag.com', 'www.christmasarchives.com', 'www.mnmidwestfoodequipment.com', 'www.etymonline.com', 'www.italymagazine.com', 'www.gallup.com', 'www.encyclopedia.com', 'books.google.com', 'www.historytoday.com', 'books.google.com', 'simplytreasures.com', 'books.google.com', 'www.christianitytoday.com', 'books.google.com', 'books.google.com', 'www.jewishworldreview.com', 'www.mnmidwestfoodequipment.com', 'www.time.com', 'www.siouxcityjournal.com', 'www.countryliving.com', 'articles.latimes.com', 'books.google.com', 'skiathosbooks.com', 'www.latimes.com', 'www.soundvision.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.gallup.com', 'www.roger-pearse.com', 'www.washingtonpost.com', 'www.nytimes.com', 'www.usatoday.com', 'www.etymonline.com', 'books.google.com', 'books.google.com', 'retailindustry.about.com', 'enduringword.com', 'books.google.com', 'www.bbc.com', 'sites.google.com', 'www.voanews.com', 'www.gardeningknowhow.com', 'www.history.com', 'books.google.com', 'www.americanstationery.com', 'books.google.com', 'books.google.com', 'www.historytoday.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.historytoday.com', 'articles.latimes.com', 'books.google.com', 'www.scribd.com', 'books.google.com', 'europe.stripes.com', 'www.etymonline.com', 'www.nbcnews.com', 'www.nbcnews.com', 'books.google.com', 'books.google.com', 'www.fashion-era.com', 'books.google.com', 'books.google.com', 'gbod-assets.s3.amazonaws.com', 'www.scmp.com', 'www.economist.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'www.forbes.com', 'books.google.com', 'www.rd.com', 'books.google.com', 'encyclopediaofukraine.com', 'www.americanstationery.com', 'www.roger-pearse.com', 'www.thehistoryofchristmas.com', 'www.christianitytoday.com', 'www.bbc.com', 'www.history.com', 'www.investopedia.com', 'womeninbusiness.about.com', 'www.etymonline.com', 'historybuff.com', 'books.google.com', 'books.google.com', 'www.enn.com', 'aclj.org', 'www.gutenberg.org', 'www.jstor.org', 'kafkadesk.org', 'www.pewforum.org', 'tertullian.org', 'www.fpchurch.org', 'www.muslimcanadiancongress.org', 'www.biblicalarchaeology.org', 'carnegiemnh.org', 'www.biblicalarchaeology.org', 'www.crivoice.org', 'www.pewforum.org', 'livius.org', 'www.catholicculture.org', 'www.belcherfoundation.org', 'www.oremus.org', 'ethiopianorthodox.org', 'www.tuc.org', 'tertullian.org', 'www.r-site.org', 'www.iwm.org', 'www.fas.org', ['harvard data science review'], ['[[grove music online', '[[oxford university press']]",6237,Require administrator access (no expiry set),191251,31 October 2001,208.235.58.xxx ,11405,14,2001-10-31,2001-10,2001
377,377,Scottish people,https://en.wikipedia.org/wiki/Scottish_people,106,0,[],[],9,20,0,26,0,0,52,0.08490566037735849,0.18867924528301888,0.24528301886792453,0.0,0.0,0.27358490566037735,0,"['www.scotlandscensus.gov', 'www.ons.gov', 'stats.gov', 'www.friendsofscotland.gov', 'www.gov', 'www.friendsofscotland.gov', 'www.gov', 'webarchive.loc.gov', 'stats.gov', 'www.gov', 'www.censusdata.abs.gov', 'www.gov', 'www.gov', 'factfinder.census.gov', 'www.scotland.gov', 'www.nrscotland.gov', 'www.scotland.gov', 'www.censusdata.abs.gov', 'stats.gov', 'www.gov', 'www.forgottenbooks.com', 'electricscotland.com', 'books.google.com', 'dictionary.com', 'answers.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.scotsman.com', 'www.heraldscotland.com', 'warsaw-life.com', 'encarta.msn.com', 'statisticalatlas.com', 'www.qldmigrationheritage.com', 'www.scotsman.com', 'www.deliciousitaly.com', 'askoxford.com', 'www.ancestralscotland.com', 'books.google.com', 'www.highbeam.com', 'www.irishtimes.com', 'www.wsj.com', 'naturemagics.com', 'books.google.com', 'electricscotland.com', 'books.google.com', 'bord-na-gaidhlig.org', 'scotland.org', 'scotland.org', 'visitscotland.org', 'scotland.org', 'www.scottishaffairs.org', 'scotland.org', 'www.aughty.org', 'strathspey.org']",34850722,Allow all users (no expiry set),80599,7 August 2004,66.185.85.80 ,3450,11,2004-08-07,2004-08,2004
378,378,Culture of Greece,https://en.wikipedia.org/wiki/Culture_of_Greece,22,1,"['10.1525/ae.1999.26.1.196', None, None]",[['american ethnologist']],0,0,0,5,0,0,16,0.0,0.0,0.22727272727272727,0.045454545454545456,0.0,0.045454545454545456,1,"['www.zeenews.com', 'dsc.discovery.com', 'm-w.com', 'www.24grammata.com', 'www.focusmm.com', ['american ethnologist']]",187260,Allow all users (no expiry set),76421,23 February 2003,195.242.150.142 ,3195,1,2003-02-23,2003-02,2003
379,379,Culture of Romania,https://en.wikipedia.org/wiki/Culture_of_Romania,7,0,[],[],0,0,0,2,0,0,5,0.0,0.0,0.2857142857142857,0.0,0.0,0.0,0,"['www.britannica.com', 'www.britannica.com']",224643,Allow all users (no expiry set),57745,10 May 2003,Bogdangiusca ,851,2,2003-05-10,2003-05,2003
380,380,Galicia (Spain),https://en.wikipedia.org/wiki/Galicia_(Spain),99,0,[],[],3,1,0,25,0,0,70,0.030303030303030304,0.010101010101010102,0.25252525252525254,0.0,0.0,0.04040404040404041,0,"['data.aad.gov', 'breathingalicia.com', 'www.parlamentodegalicia.com', 'thelatinlibrary.com', 'www.forbes.com', 'santiagoways.com', 'ccaa.elpais.com', 'www.finanzzas.com', 'www.collinsdictionary.com', 'cotizalia.com', 'www.lavanguardia.com', 'www.elespanol.com', 'www.facebook.com', 'www.xornal.com', 'www.elpais.com', 'elprogreso.galiciae.com', 'galicia-hoxe.com', 'galiciae.com', 'www.parlamentodegalicia.com', 'www.ethnologue.com', 'www.galiciaparaelmundo.com', 'www.elpais.com', 'durvate.wordpress.com', 'verne.elpais.com', 'www.cincodias.com', 'www.vieiros.com', 'weblogs.madrimasd.org', 'consellodacultura.org', 'hdi.globaldatalab.org']",12837,Allow all users (no expiry set),144530,14 November 2001,144.75.4.xxx ,3749,7,2001-11-14,2001-11,2001
381,381,Thistle,https://en.wikipedia.org/wiki/Thistle,32,6,"['10.1021/jf990326v', '10.15835/nbha4129298', None, '10.1371/journal.pone.0158117', '10.1603/022.038.0325', '10.1093/ajhp/56.12.1195', '10691655', None, '12722542', '27341588', '19508782', '10484652', None, None, None, '4920406', None, None]","[['journal of agricultural and food chemistry'], [' not bot horti agrobo '], ['j pharm belg '], ['plos one '], [' environmental entomology '], [' am j health syst pharm ']]",7,0,0,10,0,0,9,0.21875,0.0,0.3125,0.1875,0.0,0.40625,6,"['www.anitasfeast.com', 'ormiston.com', 'books.google.com', 'www.botanical.com', 'www.m-w.com', 'books.google.com', 'www.luontoportti.com', 'books.google.com', 'visitscotland.com', 'books.google.com', 'xerces.org', 'en.wikisource.org', 'mooc.tela-botanica.org', 'tolweb.org', 'www.butterfly-conservation.org', 'www.hear.org', 'www.conservationgrade.org', ['journal of agricultural and food chemistry'], [' not bot horti agrobo '], ['j pharm belg '], ['plos one '], [' environmental entomology '], [' am j health syst pharm ']]",2193890,Allow all users (no expiry set),25341,8 July 2005,MPF ,572,1,2005-07-08,2005-07,2005
382,382,Medellín,https://en.wikipedia.org/wiki/Medell%C3%ADn,97,1,"['10.2307/3105262', None, None]","[['the johns hopkins university press and the [[society for the history of technology', '[[technology and culture']]",19,13,0,37,0,0,28,0.1958762886597938,0.13402061855670103,0.38144329896907214,0.010309278350515464,0.0,0.3402061855670103,1,"['www.dane.gov', 'www.dane.gov', 'www.ideam.gov', 'www.dane.gov', 'www.dane.gov', 'www.dane.gov', 'metroplus.gov', 'www.ideam.gov', 'www.dane.gov', 'www.dane.gov', 'www.ideam.gov', 'www.rosario.gov', 'www.medellin.gov', 'rankings.americaeconomia.com', 'www.lanacion.com', 'www.argos.com', 'eltiempo.com', 'www.americalate.com', 'www.coltejer.com', 'online.wsj.com', 'elcolombiano.com', 'emporis.com', 'www.ada-aero.com', 'abc.com', 'moovitapp.com', 'eltiempo.com', 'www.wca.com', 'americalate.com', 'books.google.com', 'www.straitstimes.com', 'www.flightglobal.com', 'www.caracol.com', 'www.huffingtonpost.com', 'eltiempo.com', 'caracol.com', 'www.metrocuadrado.com', 'content.time.com', 'www.elcolombiano.com', 'www.proexport.com', 'albeiror24.wordpress.com', 'pbfernandobotero.blogspot.com', 'www.leekuanyewworldcityprize.com', 'www.tuneldeoccidente.com', 'suleasing-intl.com', 'sostenibilidad.semana.com', 'books.google.com', 'travel.nationalgeographic.com', 'moovitapp.com', 'www.touringmedellin.com', 'www.llworldtour.com', 'www.reddebibliotecas.org', 'ciudaddonbosco.org', 'www.sister-cities.org', 'socearq.org', 'creativetourismnetwork.org', 'creativecommons.org', 'igarape.org', 'www.itdp.org', 'www.unhabitat.org', 'www.cipcol.org', 'www.gatesfoundation.org', 'brtdata.org', 'www.camaramed.org', 'www.odi.org', 'rightlivelihood.org', 'www.globalurban.org', 'seguridadjusticiaypaz.org', 'www.olympic.org', '54pesos.org', ['the johns hopkins university press and the [[society for the history of technology', '[[technology and culture']]",340197,Allow all users (no expiry set),134099,13 October 2003,Jaleho ,3235,6,2003-10-13,2003-10,2003
383,383,Culture of Germany,https://en.wikipedia.org/wiki/Culture_of_Germany,84,1,"[None, 'kmeigen.kmpresse_1408435283&start=0&anzahl=10&channel=kmeigen&language=e&archiv=', None]",[['gamescom press center']],10,1,0,29,0,1,42,0.11904761904761904,0.011904761904761904,0.34523809523809523,0.011904761904761904,0.0,0.14285714285714285,1,"['www.centennialofflight.gov', 'www.bbc.com', 'www.gaycitynews.com', 'www.news24.com', 'www.gaycitynews.com', 'www.nationmaster.com', 'encarta.msn.com', 'www.filmbug.com', 'www.britannica.com', 'archive.wired.com', 'in.reuters.com', 'economictimes.indiatimes.com', 'dw.com', 'www.epemag.com', 'gizmodo.com', 'www.pyeongchang2018.com', 'cooking.nytimes.com', 'www.tourism-review.com', 'www.german-way.com', 'www.nationmaster.com', 'www.gfk.com', 'www.german-way.com', 'royalunibrew.com', 'www.history.com', 'dw.com', 'rio2016.com', 'books.google.com', 'www.howtogermany.com', 'www.imdb.com', 'de.statista.com', 'www.jewishvirtuallibrary.org', 'www.fiapf.org', 'worldpublicopinion.org', 'www.germanhistorydocs.ghi-dc.org', 'worldpublicopinion.org', 'www.alumniportal-deutschland.org', 'germanfoods.org', 'www.worldheritagesite.org', 'www.org', 'www.alumniportal-deutschland.org', ['gamescom press center']]",1195868,Allow all users (no expiry set),62654,22 November 2004,Sextus~enwiki ,1556,0,2004-11-22,2004-11,2004
384,384,Rize Province,https://en.wikipedia.org/wiki/Rize_Province,24,0,[],[],2,0,0,9,0,0,13,0.08333333333333333,0.0,0.375,0.0,0.0,0.08333333333333333,0,"['www.encyclopedia.com', 'www.karalahana.com', 'www.nytimes.com', 'www.karalahana.com', 'www.karalahana.com', 'www.weatherbase.com', 'www.dailysabah.com', 'www.dailysabah.com', 'karalahana.com', 'www.iranicaonline.org', 'dergipark.org']",886778,Allow all users (no expiry set),22875,8 August 2004,Avnionur ,339,0,2004-08-08,2004-08,2004
385,385,Odia people,https://en.wikipedia.org/wiki/Odia_people,16,0,[],[],0,2,0,13,0,0,1,0.0,0.125,0.8125,0.0,0.0,0.125,0,"['www.censusindia.gov', 'www.censusindia.gov', 'books.google.com', 'www.dailypioneer.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'thenewleam.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehindu.com', 'www.ethnologue.com', 'books.google.com', 'odishanewsinsight.com', 'telanganatoday.com']",5210850,Require administrator access (no expiry set),27670,19 May 2006,Afghan Historian ,1126,2,2006-05-19,2006-05,2006
386,386,Dolphin,https://en.wikipedia.org/wiki/Dolphin,230,35,"['10.1098/rsbl.2018.0314', '10.1213/01.ane.0000250369.33700.eb', '10.3389/fphys.2020.604018', '10.1007/s00359-013-0817-7', '10.1002/ar.20407', '10.1111/j.1751-0813.2011.00849.x', '10.1038/nature06343', '10.1002/ar.20528', '10.1017/s0025315407054215', '10.1073/pnas.1108927108', '10.1016/j.meegid.2011.08.018', '10.1007/978-3-642-69554-4_17', '10.1073/pnas.0409518102', '10.1037/0735-7036.114.1.98', '10.1163/1568539053627712', '10.1126/science.aat4220', '10.3819/ccbr.2008.30003', '10.1177/030098586900600307', '10.1016/j.neuroscience.2006.04.084', '10.1016/j.icesjms.2005.06.012', '10.1242/jeb.203.14.2125', '10.1111/j.1439-0442.2005.00693.x', '10.1093/icb/42.5.1071', '10.1017/s0025315407055233', '10.1136/bmj.331.7527.1231', '10.1002/ar.20529', '10.1037/0735-7036.122.3.305', '10.1146/annurev.ecolsys.33.020602.095426', '10.1007/s10914-011-9184-8', '10.1006/ccog.1995.1026', '10.1016/j.tics.2005.06.008', '10.1016/s1095-6433(00)00182-3', '10.1136/bmj.331.7529.1407', '10.2752/089279307x224782', '30185606', '17179314', '33329056', '23649908', '17441195', '22008125', '18097400', '17516434', None, '21873217', '21888991', None, '15677331', '10739315', None, '30679341', None, '5817449', '16797136', None, '10862725', '15737178', '21680390', None, '16308382', '17516421', '18729659', None, None, '8521259', '16002323', '10936758', '16339258', None, '6170752', None, '7732665', None, None, None, None, None, None, '3167538', None, None, '547867', None, None, None, None, None, None, None, None, None, None, None, '1289317', None, None, None, None, None, None, None, '1309662', None]","[[' [[biol lett.'], ['anesthesia '], ['[[frontiers in physiology'], ['journal of comparative physiology'], ['the anatomical record '], [' australian veterinary journal '], ['nature '], ['the anatomical record '], ['journal of the marine biological association of the uk'], ['pnas '], [' infection'], ['experimental brain research'], ['proceedings of the national academy of sciences '], ['journal of comparative psychology '], ['behaviour'], ['science'], ['comparative cognition '], ['veterinary pathology'], ['neuroscience '], [' ices journal of marine science'], ['journal of experimental biology '], [' journal of veterinary medicine'], ['integrative and comparative biology '], [' journal of the marine biological association of the uk'], ['bmj '], ['anatomical record '], ['journal of comparative psychology'], ['annual review of ecology and systematics '], ['journal of mammalian evolution '], ['consciousness and cognition'], ['trends cogn sci '], [' comparative biochemistry and physiology. part a'], [' bmj'], ['anthrozoös ']]",26,3,0,54,0,2,110,0.11304347826086956,0.013043478260869565,0.23478260869565218,0.15217391304347827,0.0,0.2782608695652174,34,"['india.gov', 'swfsc.noaa.gov', 'www.nmfs.noaa.gov', 'atlantisthepalm.com', 'yellowmagpie.com', 'www.nytimes.com', 'www.adelaidenow.com', 'www.cbsnews.com', 'www.newscientist.com', 'asiancorrespondent.com', 'www.youtube.com', 'wordnik.com', 'www.youtube.com', 'www.cnn.com', 'www.seeker.com', 'www.nytimes.com', 'www.hakaimagazine.com', 'www.nytimes.com', 'www.trustedpartner.com', 'livescience.com', 'dolphinmovie.com', 'articles.orlandosentinel.com', 'www.youtube.com', 'www.reuters.com', 'dictionary.reference.com', 'news.discovery.com', 'www.atuna.com', 'www.juneauempire.com', 'dw.com', 'www.news.com', 'www.watoday.com', 'dolphinsafari.com', 'www.wired.com', 'news.nationalgeographic.com', 'www.sciencedaily.com', 'www.healthline.com', 'www.livescience.com', 'news.nationalgeographic.com', 'blogs.scientificamerican.com', 'cookpad.com', 'www.vice.com', 'www.huffingtonpost.com', 'www.cnn.com', 'www.nationalgeographic.com', 'www.dolphindock.com', 'www.bbc.com', 'www.livescience.com', 'science-frontiers.com', 'www.txtwriter.com', 'today.msnbc.msn.com', 'news.nationalgeographic.com', 'blogs.discovermagazine.com', 'animals.mom.com', 'dictionary.com', 'www.nytimes.com', 'www.irishcentral.com', 'cracked.com', 'nmmpfoundation.org', 'acsonline.org', 'www.pnas.org', 'fishingnj.org', 'animalquestions.org', 'www.whalefacts.org', 'www.pbs.org', 'marineconservation.org', 'www.afd.org', 'www.elasmo-research.org', 'us.whales.org', 'islandheritage.org', 'www.tmmsn.org', 'phys.org', 'seaworld.org', 'portals.iucn.org', 'www.hsi.org', 'www.fishbase.org', 'www.humanesociety.org', 'whalesalive.org', 'mbe.oxfordjournals.org', 'sharkangels.org', 'hsi.org', 'acsonline.org', 'marinebio.org', 'www.robins-island.org', [' [[biol lett.'], ['anesthesia '], ['[[frontiers in physiology'], ['journal of comparative physiology'], ['the anatomical record '], [' australian veterinary journal '], ['nature '], ['the anatomical record '], ['journal of the marine biological association of the uk'], ['pnas '], [' infection'], ['experimental brain research'], ['proceedings of the national academy of sciences '], ['journal of comparative psychology '], ['behaviour'], ['science'], ['comparative cognition '], ['veterinary pathology'], ['neuroscience '], [' ices journal of marine science'], ['journal of experimental biology '], [' journal of veterinary medicine'], ['integrative and comparative biology '], [' journal of the marine biological association of the uk'], ['bmj '], ['anatomical record '], ['journal of comparative psychology'], ['annual review of ecology and systematics '], ['journal of mammalian evolution '], ['consciousness and cognition'], ['trends cogn sci '], [' comparative biochemistry and physiology. part a'], [' bmj'], ['anthrozoös ']]",9061,Require administrator access (no expiry set),124958,1 January 2002,Di Stroppo ,3952,2,2002-01-01,2002-01,2002
387,387,Djibouti,https://en.wikipedia.org/wiki/Djibouti,153,6,"['10.1525/ae.1975.2.4.02a00030', '10.3406/ethio.1987.931', '10.3406/cea.1968.3123', '10.1029/96jb01185', None, None, None, None, None, None, None, None]","[['american ethnologist '], ['annales d'], ['cahiers d'], ['journal of geophysical research']]",27,6,0,58,0,0,56,0.17647058823529413,0.0392156862745098,0.3790849673202614,0.0392156862745098,0.0,0.2549019607843137,4,"['www.cia.gov', 'www.cia.gov', 'www.cia.gov', 'lcweb2.loc.gov', 'eastafrica.usaid.gov', 'www.cia.gov', 'allafrica.com', 'www.awdalpress.com', 'www.nytimes.com', 'theculturetrip.com', 'books.google.com', 'www.cbsnews.com', 'ethiosports.com', 'image.prntsacr.com', 'historyorb.com', 'books.google.com', 'basementgeographer.com', 'lntreasures.com', 'www.worldatlas.com', 'books.google.com', 'www.scmp.com', 'www.google.com', 'www.google.com', 'www.middle-east-online.com', 'www.africanews.com', 'www.google.com', 'www.reuters.com', 'www.google.com', 'books.google.com', 'allafrica.com', 'www.eiu.com', 'books.google.com', 'www.google.com', 'www.weatherbase.com', 'www.businessdailyafrica.com', 'books.google.com', 'books.google.com', '2rep.legion-etrangere.com', 'books.google.com', 'books.google.com', 'goobjoog.com', 'www.google.com', 'www.britannica.com', 'www.google.com', 'www.google.com', 'defaakto.com', 'bloomberg.com', 'www.google.com', 'www.euromoneycountryrisk.com', 'www.cnbc.com', 'books.google.com', 'books.google.com', 'www.ethnologue.com', 'steelguru.com', 'sabahionline.com', 'books.google.com', 'books.google.com', 'www.onceinalifetimejourney.com', 'www.oxfordbusinessgroup.com', 'www.nytimes.com', 'www.google.com', 'www.awdalpress.com', 'www.oxfordreference.com', 'books.google.com', 'djibouti.frontafrique.org', 'www.irinnews.org', 'www.aaeafrica.org', 'www.unfpa.org', 'www.freedomhouse.org', 'www.jstor.org', 'cinematreasures.org', 'hdr.undp.org', 'www.wfp.org', 'catholic-hierarchy.org', 'www.un.org', 'www.nationsonline.org', 'www.imf.org', 'djibouti.frontafrique.org', 'somavires.org', 'whc.unesco.org', 'www.constituteproject.org', 'www.infodev.org', 'geonames.org', 'www.pewforum.org', 'www.chathamhouse.org', 'www.irinnews.org', 'pewforum.org', 'documents.worldbank.org', 'www.irinnews.org', 'www.refworld.org', 'unhcr.org', ['american ethnologist '], ['annales d'], ['cahiers d'], ['journal of geophysical research']]",17207794,Require administrator access (no expiry set),130003,26 April 2001,KoyaanisQatsi ,6069,1,2001-04-26,2001-04,2001
388,388,Mallorca,https://en.wikipedia.org/wiki/Mallorca,93,5,"['10.1038/s41559-020-1102-0', '10.1177/09596836211060491', '10.1080/01434632.2014.979832', '10.1007/s10963-008-9010-2', '10.24965/da.v0i3.10371', '32094539', None, None, None, None, '7080320', None, None, None, None]","[['nature ecology '], ['the holocene'], ['journal of multilingual and multicultural development'], ['journal of world prehistory'], ['documentación administrativa', '[[instituto nacional de administración pública']]",3,1,0,38,0,1,45,0.03225806451612903,0.010752688172043012,0.40860215053763443,0.053763440860215055,0.0,0.0967741935483871,5,"['www.me.gov', 'elpais.com', 'www.abc-mallorca.com', 'www.majorca.com', 'www.alcudia-boat-rental.com', 'www.majorcanvillas.com', 'www.collinsdictionary.com', 'www.vipealo.com', 'books.google.com', 'allthatsinteresting.com', 'elpais.com', 'mallorcaincognita.com', 'www.contemporarybalears.com', 'www.elcultural.com', 'answers.com', 'www.ludwig-salvator.com', 'mallorcaincognita.com', 'politica.elpais.com', 'dw.com', 'www.northsouthguides.com', 'www.papelesdesonarmadans.com', 'www.helencummins.com', 'www.lavanguardia.com', 'www.abc-mallorca.com', 'es.ripleybelieves.com', 'worldatlas.com', 'politica.elpais.com', 'www.alcudia-boat-rental.com', 'www.dw.com', 'www.weather-atlas.com', 'www.seemallorca.com', 'www.mallorcaaventura.com', 'www.cntraveler.com', 'www.lonelyplanet.com', 'talksport.com', 'www.majorcadailybulletin.com', 'www.typicallyspanish.com', 'www.myguidemallorca.com', 'cafebabel.com', 'whc.unesco.org', 'om.ciheam.org', 'seatemperature.org', ['nature ecology '], ['the holocene'], ['journal of multilingual and multicultural development'], ['journal of world prehistory'], ['documentación administrativa', '[[instituto nacional de administración pública']]",59310,Allow all users (no expiry set),77029,24 June 2002,Jeronimo ,3010,2,2002-06-24,2002-06,2002
389,389,Bengal,https://en.wikipedia.org/wiki/Bengal,158,4,"['10.1109/mwsym.1997.602854', '10.2307/2642858', '10.2307/3454378', '10.1007/bf00175563', None, None, '10811564', None, None, None, '1638054', None]","[['ieee '], ['asian survey '], ['[[environmental health perspectives'], ['water']]",24,17,0,74,0,1,38,0.1518987341772152,0.10759493670886076,0.46835443037974683,0.02531645569620253,0.0,0.2848101265822785,4,"['censusindia.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'www.mea.gov', 'www.censusindia.gov', 'www.cia.gov', 'www.censusindia.gov', 'bdlaws.minlaw.gov', 'www.censusindia.gov', 'memory.loc.gov', 'www.censusindia.gov', 'www.bbs.gov', 'www.vigyanprasar.gov', 'censusindia.gov', 'www.censusindia.gov', 'censusindia.gov', 'www.censusindia.gov', 'www.britannica.com', 'indianmirror.com', 'books.google.com', 'books.google.com', 'www.ethnologue.com', 'books.google.com', 'www.nytimes.com', 'en.oxforddictionaries.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.bbc.com', 'global.britannica.com', 'www.wbtourism.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'thediplomat.com', 'books.google.com', 'books.google.com', 'books.google.com', 'storyofpakistan.com', 'www.etymonline.com', 'books.google.com', 'books.google.com', 'www.asansolmunicipalcorporation.com', 'link.galegroup.com', 'books.google.com', 'wanderinggaia.com', 'storyofpakistan.com', 'books.google.com', 'archive.dhakatribune.com', 'books.google.com', 'importantindia.com', 'books.google.com', 'www.livemint.com', 'books.google.com', 'www.britannica.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'books.google.com', 'news.xinhuanet.com', 'www.hinduonnet.com', 'nation.com', 'books.google.com', 'books.google.com', 'copenhagenconsensus.com', 'www.thaindian.com', 'books.google.com', 'books.google.com', 'www.reuters.com', 'newagebd.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'factsanddetails.com', 'www.bbc.com', 'books.google.com', 'www.livemint.com', 'books.google.com', 'books.google.com', 'articles.economictimes.indiatimes.com', 'bengalonline.sitemarvel.com', 'books.google.com', 'books.google.com', 'books.google.com', 'en.banglapedia.org', 'en.banglapedia.org', 'www.sciencehistory.org', 'metmuseum.org', 'cri.org', 'akdn.org', 'worldviewcities.org', 'www.org', 'en.banglapedia.org', 'en.banglapedia.org', 'worldviewcities.org', 'www.unicef.org', 'www.yhaindia.org', 'en.banglapedia.org', 'en.banglapedia.org', 'www.rbi.org', 'en.banglapedia.org', 'en.banglapedia.org', 'en.banglapedia.org', 'en.banglapedia.org', 'www.saarc-sec.org', 'www.worldcat.org', 'govdocs.aquake.org', 'en.banglapedia.org', ['ieee '], ['asian survey '], ['[[environmental health perspectives'], ['water']]",4862,"Require autoconfirmed or confirmed access (18:26, 29 June 2023)",134218,22 December 2001,Hagedis ,3241,6,2001-12-22,2001-12,2001
390,390,Mycenaean Greece,https://en.wikipedia.org/wiki/Mycenaean_Greece,353,24,"['10.2307/504929', '10.1007/bf00140587', '10.1111/1468-0092.00084', '10.2307/148143', '10.2307/506802', '10.2307/504928', '10.1017/s006824540001409x', '10.1353/are.2015.0007', '10.2307/505489', '10.1111/j.1468-0092.1996.tb00087.x', '10.1017/ccol9780521814447.011', '10.1038/nature23310', '10.1006/jasc.1999.0431', '10.11588/diglit.811', '10.3406/ahess.1982.282879', 'abs/10.1002/jqs.3314', '10.1017/s0003598x00041740', '10.2143/bib.101.3.3288731', '10.2972/hesperia.86.4.0583', '10.1111/j.2041-5370.1999.tb00480.x', '10.1017/s0003598x00040187', '10.1080/00497878.1981.9978529', '10.11141/ia.56.9', None, None, None, None, None, None, None, None, None, None, None, '28783727', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, '5565772', None, None, None, None, None, None, None, None, None, None, None]","[['american journal of archaeology'], ['climatic change'], ['oxford journal of archaeology'], ['hesperia'], ['[[american journal of archaeology'], ['american journal of archaeology'], ['annual of the british school at athens'], ['arethusa'], ['american journal of archaeology'], ['oxford journal of archaeology'], ['cambridge university press'], ['nature'], ['journal of archaeological science'], ['macmillan'], ['annales. histoire'], ['journal of quaternary science'], ['antiquity'], ['biblica '], ['hesperia'], ['bulletin of the institute of classical studies'], ['antiquity'], ['women'], ['internet archaeology']]",7,0,0,70,0,0,252,0.019830028328611898,0.0,0.19830028328611898,0.0679886685552408,0.0,0.08781869688385269,23,"['books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.salimbeti.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.livescience.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.cbsnews.com', 'www.britannica.com', 'www.livescience.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'submissions.e-a-a.org', 'www.sciencemag.org', 'www.sbl-site.org', 'phys.org', 'www.worldhistory.org', 'submissions.e-a-a.org', 'www.metmuseum.org', ['american journal of archaeology'], ['climatic change'], ['oxford journal of archaeology'], ['hesperia'], ['[[american journal of archaeology'], ['american journal of archaeology'], ['annual of the british school at athens'], ['arethusa'], ['american journal of archaeology'], ['oxford journal of archaeology'], ['cambridge university press'], ['nature'], ['journal of archaeological science'], ['macmillan'], ['annales. histoire'], ['journal of quaternary science'], ['antiquity'], ['biblica '], ['hesperia'], ['bulletin of the institute of classical studies'], ['antiquity'], ['women'], ['internet archaeology']]",565602,Allow all users (no expiry set),135638,31 March 2004,Adam Carr ,2465,6,2004-03-31,2004-03,2004
391,391,Yunnan,https://en.wikipedia.org/wiki/Yunnan,100,8,"['10.1007/s10722-021-01309-y', '10.3406/adh.1982.1543', '10.1016/j.pld.2020.07.006', '10.1023/b:bioc.0000011728.46362.3c', None, '10.3897/zookeys.864.26689', '10.1007/s10531-013-0579-0', '10.1007/s10764-009-9360-3', None, None, None, None, '23913883', '31363346', None, '19644553', None, None, None, None, None, '6656784', None, '2715875']","[['genetic resources and crop evolution '], ['annales de démographie historique '], ['plant diversity '], ['biodiversity '], [' dong wu xue yan jiu '], ['zookeys ', 'pensoft publishers '], ['biodiversity and conservation'], [' international journal of primatology']]",11,15,0,19,0,1,46,0.11,0.15,0.19,0.08,0.0,0.34,8,"['stats.yn.gov', 'www.stats.gov', 'www.nmc.gov', 'www.stats.gov', 'data.stats.gov', 'www.sztj.gov', 'english.mofcom.gov', 'www.sztj.gov', 'data.stats.gov', 'www.stats.gov', 'www.stats.gov', 'www.stats.gov', 'www.stats.gov', 'files2.mca.gov', 'www.stats.gov', 'books.google.com', 'www.ttgmice.com', 'books.google.com', 'www.kmgairport.com', 'yn.cppiae.com', 'thechinaperspective.com', 'books.google.com', 'books.google.com', 'www.thecultureconcept.com', 'www.nytimes.com', 'books.google.com', 'windrug.com', 'books.google.com', 'www.history.com', 'english.people.com', 'news.xinhuanet.com', 'www.reuters.com', 'books.google.com', 'urbandwellerscoffee.com', 'globaldatalab.org', 'alertnet.org', 'whc.unesco.org', 'www.usp.org', 'portal.unesco.org', 'www.kunming.org', 'baylor-ir.tdl.org', 'www.gutenberg-e.org', 'www.china.org', 'the-leaf.org', 'www.wdl.org', ['genetic resources and crop evolution '], ['annales de démographie historique '], ['plant diversity '], ['biodiversity '], [' dong wu xue yan jiu '], ['zookeys ', 'pensoft publishers '], ['biodiversity and conservation'], [' international journal of primatology']]",166410,Allow all users (no expiry set),124969,7 January 2003,Olivier ,1780,4,2003-01-07,2003-01,2003
392,392,Culture of Iraq,https://en.wikipedia.org/wiki/Culture_of_Iraq,18,3,"['10.5622/illinois/9780252041280.003.0005', '10.4324/9781315474618-6', None, None, None, None]","[['university of illinois press'], ['routledge']]",3,0,0,7,0,0,5,0.16666666666666666,0.0,0.3888888888888889,0.16666666666666666,0.0,0.3333333333333333,2,"['books.google.com', 'www.xinhuanet.com', 'books.google.com', 'www.britannica.com', 'www.pilotguides.com', 'insidearabia.com', 'www.thingsasian.com', 'www.worldcat.org', 'www.worldcat.org', 'www.worldcat.org', ['university of illinois press'], ['routledge']]",176531,Allow all users (no expiry set),25622,30 January 2003,64.12.96.13 ,749,2,2003-01-30,2003-01,2003
393,393,Guatemala,https://en.wikipedia.org/wiki/Guatemala,218,4,"['10.1017/s000316150008843x', '10.1215/01636545-1994-58-35', '10.1177/0094582x9902600207', '10.1038/s41467-020-19493-3', None, None, None, '33293507', None, None, None, '7723057']","[['the americas', 'academy of american franciscan history'], ['radical history review'], ['latin american perspectives'], ['nature communications']]",46,4,0,85,0,1,79,0.21100917431192662,0.01834862385321101,0.38990825688073394,0.01834862385321101,0.0,0.24770642201834864,4,"['www.justice.gov', 'www.cia.gov', 'pdf.usaid.gov', 'www.state.gov', 'www1.folha.uol.com', 'www.haaretz.com', 'm.elperiodico.com', 'www.reuters.com', 'books.google.com', 'books.google.com', 'www.s21.com', 'www.nytimes.com', 'www.prensalibre.com', 'www.nytimes.com', 'www.docstoc.com', 'www.nytimes.com', 'weather.com', 'bgr.com', 'www.thearda.com', 'www.bbc.com', 'bbcnews.com', 'www.prensalibre.com', 'www.bbc.com', 'latinartmuseum.com', 'www.prensalibre.com', 'www.prensalibre.com', 'www.bbc.com', 'books.google.com', 'servicios.prensalibre.com', 'www.scribd.com', 'www.history.com', 'www.elperiodico.com', 'www.fivb.com', 'www.s21.com', 'www.reuters.com', 'books.google.com', 'www.washingtonpost.com', 'dw.com', 'www.cervantesvirtual.com', 'msn.com', 'books.google.com', 'yahoo.com', 'books.google.com', 'www.newsweek.com', 'latinartmuseum.com', 'books.google.com', 'books.google.com', 'time.com', 'www.deguate.com', 'datosmacro.expansion.com', 'www.nytimes.com', 'www.nytimes.com', 'books.google.com', 'elperiodico.com', 'www.guatemalago.com', 'www.bbc.com', 'magazine.mining.com', 'books.google.com', 'www.authenticmaya.com', 'naranetacrossing.wordpress.com', 'www.routledge.com', 'rainforestcentralamerica.wordpress.com', 'elperiodico.com', 'www.newsweek.com', 'books.google.com', 'books.google.com', 'www.christianitytoday.com', 'olodonation.com', 'www.prensalibre.com', 'www.bbc.com', 'www.prensalibre.com', 'www.nytimes.com', 'books.google.com', 'www.plazapublica.com', 'www.guatevision.com', 'noticias.emisorasunidas.com', 'evangelicalfocus.com', 'www.ancientfaith.com', 'www.washingtonpost.com', 'ldschurchtemples.com', 'www.businessinsider.com', 'datosmacro.expansion.com', 'elperiodico.com', 'www.nytimes.com', 'prensalibre.com', 'books.google.com', 'noticias.emisorasunidas.com', 'www.prensalibre.com', 'www.nationalgeographic.com', 'bibliolore.org', 'www.unesco.org', 'shr.aaas.org', 'www.iucn.org', 'www.afehc-historia-centroamericana.org', 'data.worldbank.org', 'www.insightcrime.org', 'commons.wikimedia.org', 'www.migrationdrc.org', 'www.cicig.org', 'www.ppu.org', 'www.democracynow.org', 'migrationinformation.org', 'www.goarchmexico.org', 'www.sciencenews.org', 'www.albedrio.org', 'churchofjesuschrist.org', 'www.biodiversityhotspots.org', 'www.asil.org', 'www.albedrio.org', 'www.insightcrime.org', 'stats.uis.unesco.org', 'catalog.hathitrust.org', 'hdr.undp.org', 'cmiguate.org', 'hdr.undp.org', 'hdr.undp.org', 'iucn.org', 'www.refworld.org', 'www.famsi.org', 'nacla.org', 'www.focolare.org', 'www.insightcrime.org', 'data.worldbank.org', 'www.albedrio.org', 'web.worldbank.org', 'imf.org', 'churchofjesuschristtemples.org', 'web.amnesty.org', 'esa.un.org', 'ccidinc.org', 'treaties.un.org', 'hdr.undp.org', 'documents.worldbank.org', 'econ.worldbank.org', 'web.amnesty.org', ['the americas', 'academy of american franciscan history'], ['radical history review'], ['latin american perspectives'], ['nature communications']]",17238567,Require administrator access (no expiry set),184724,10 September 2001,Koyaanis Qatsi ,10438,17,2001-09-10,2001-09,2001
394,394,Prato,https://en.wikipedia.org/wiki/Prato,15,0,[],[],0,0,0,6,0,0,9,0.0,0.0,0.4,0.0,0.0,0.0,0,"['www.nytimes.com', 'www.com', 'articles.chicagotribune.com', 'www.textileworld.com', 'adribarrcrocetti.com', 'www.com']",1821975,Allow all users (no expiry set),28260,30 April 2005,Dryazan ,676,4,2005-04-30,2005-04,2005
395,395,Culture of Belgium,https://en.wikipedia.org/wiki/Culture_of_Belgium,37,0,[],[],5,0,0,22,0,0,10,0.13513513513513514,0.0,0.5945945945945946,0.0,0.0,0.13513513513513514,0,"['www.visitbelgium.com', 'articles.chicagotribune.com', 'www.inbev.com', 'www.epicurious.com', 'www.globalgourmet.com', 'wwar.com', 'www.senses-artnouveau.com', 'wwar.com', 'www.senses-artnouveau.com', 'fashionworlds.blogspot.com', 'www.belgianexperts.com', 'wwar.com', 'www.belgianexperts.com', 'wwar.com', 'www.britannica.com', 'www.epicurious.com', 'www.globalgourmet.com', 'www.globalpost.com', 'www.filmbirth.com', 'houbi.com', 'www1.uol.com', 'www.filmbirth.com', 'whc.unesco.org', 'www.metmuseum.org', 'www.metmuseum.org', 'www.unesco.org', 'www.metmuseum.org']",143432,Allow all users (no expiry set),32343,3 November 2002,12.233.64.10 ,574,9,2002-11-03,2002-11,2002
396,396,Culture of Wales,https://en.wikipedia.org/wiki/Culture_of_Wales,143,0,[],[],13,3,0,37,0,4,86,0.09090909090909091,0.02097902097902098,0.25874125874125875,0.0,0.0,0.11188811188811189,0,"['cadw.gov', 'www.rcahmw.gov', 'www.wrexham.gov', 'www.visual-arts-cork.com', 'www.welshpremier.com', 'www.economist.com', 'books.google.com', 'books.google.com', 'www.mtv.com', 'books.google.com', 'books.google.com', 'uk.com', 'books.google.com', 'books.google.com', 'books.google.com', 'photography.nationalgeographic.com', 'llantrisantchoir.com', 'allaboutartschools.com', 'www.microsofttranslator.com', 'louisekosman.com', 'www.canugwerin.com', 'books.google.com', 'www.fifa.com', 'www.royalalberthall.com', 'cardiffmalechoir.wordpress.com', 'www.historytoday.com', 'literati.credoreference.com', 'www.bbc.com', 'literati.credoreference.com', 'literati.credoreference.com', 'books.google.com', 'books.google.com', 'www.glamorgancricket.com', 'www.officialcharts.com', 'books.google.com', 'www.itv.com', 'allaboutartschools.com', 'www.officialcharts.com', 'books.google.com', 'www.microsofttranslator.com', 'imagingthebible.llgc.org', 'cerdd-dant.org', 'welshicons.org', 'www.tate.org', 'www.welshsports.org', 'herefordcathedral.org', 'www.bwwsociety.org', 'www.rcaconwy.org', 'pendyrus.org', 'www.educationengland.org', 'www.wno.org', 'www.jonathanedwards.org', 'www.cricketwales.org']",173451,Allow all users (no expiry set),71031,23 January 2003,GrahamN ,773,3,2003-01-23,2003-01,2003
397,397,Trieste,https://en.wikipedia.org/wiki/Trieste,127,1,"['10.2307/497017', None, None]",[['american journal of archaeology']],7,1,0,21,0,0,97,0.05511811023622047,0.007874015748031496,0.16535433070866143,0.007874015748031496,0.0,0.07086614173228346,1,"['www.foia.cia.gov', 'www.numbeo.com', 'www.aznations.com', 'moovitapp.com', 'www.triestecoffeecluster.com', 'www.kozina.com', 'books.google.com', 'moovitapp.com', 'books.google.com', 'books.google.com', 'www.collinsdictionary.com', 'books.google.com', 'monocle.com', 'triestetimes.com', 'www.lonelyplanet.com', 'italicsmag.com', 'www.vogue.com', 'www.collinsdictionary.com', 'books.google.com', 'eu.usatoday.com', 'www.tal-oil.com', 'www.com', 'www.deathcamps.org', 'maps.bpl.org', 'www.nzetc.org', 'www.stazionerogers.org', 'www.nuovolitorale.org', 'www.sciencefictionfestival.org', 'en.climate-data.org', ['american journal of archaeology']]",56092,Allow all users (no expiry set),110184,11 June 2002,Peterlin~enwiki ,2911,6,2002-06-11,2002-06,2002
398,398,Uyghurs,https://en.wikipedia.org/wiki/Uyghurs,379,33,"['10.1080/02634939108400758', '10.1002/elps.201800019', '10.1093/oxfordjournals.cjilaw.a000538', '10.1093/molbev/msh238', '10.1017/s0021911812000629', '10.1093/molbev/msx177', '10.1163/146481705793646892', '10.2307/1796091', '10.1016/j.ajhg.2008.08.001', '10.1080/00963402.2020.1846417', '10.1093/rsq/hdi0223', '10.1080/02634937.2012.671993', '10.1080/03071847.2020.1723284', '10.1017/s1468109915000377', '10.5038/1911-9933.15.1.1834', '10.1080/13602001003650648', '10.1002/jmv.24240', '10.1080/13602004.2012.744172', '10.1017/s0305741010000275', '10.1534/genetics.105.054270', '10.1080/0048721x.2021.1865616', '10.1016/j.ajhg.2009.10.024', '10.2753/ppc1075-8216540304', '10.1038/srep19998', '10.1080/00343404.2019.1575506', '10.1016/j.ajhg.2008.01.017', '10.1080/03068374.2019.1672433', '10.1080/10670564.2013.766383', '10.1515/opth-2015-0016', '10.1080/14631369.2010.510877', '10.1186/1471-2156-14-100', '10.1017/s0041977x00013811', None, '29869338', None, '15317881', None, '28595347', None, None, '18760393', None, None, None, None, None, None, None, '26081269', None, None, '16489223', None, '20004770', None, '26842947', None, '18355773', None, None, None, None, '24103151', None, None, None, None, None, None, None, None, None, '2556439', None, None, None, None, None, None, None, '5033003', None, None, '1456369', None, '2790568', None, '4740765', None, '2427216', None, None, None, None, '3852047', None]","[['central asian survey '], ['electrophoresis'], ['chinese journal of international law '], ['mol biol evol '], ['the journal of asian studies '], ['molecular biology and evolution'], [' inner asia ', 'brill '], ['the geographical journal'], ['americanjournal of human genetics '], ['[[bulletin of the atomic scientists'], ['refugee survey quarterly '], ['central asian survey '], ['[[rusi journal'], ['japanese journal of political science '], ['genocide studies and prevention'], ['journal of muslim minority affairs '], ['journal of medical virology '], ['journal of muslim minority affairs '], [' china quarterly '], ['genetics '], ['religion'], ['american journal of human genetics'], ['problems of post-communism '], ['scientific reports'], ['regional studies '], ['american journal of human genetics'], ['[[asian affairs'], ['journal of contemporary china '], ['open theology'], ['asian ethnicity '], ['bmc genetics'], ['bulletin of the school of oriental and african studies', 'cambridge university press on behalf of school of oriental and african studies']]",30,10,0,203,0,9,94,0.079155672823219,0.026385224274406333,0.5356200527704486,0.0870712401055409,0.0,0.19261213720316622,32,"['www.stats.gov', 'www.mfa.gov', '2001.ukrcensus.gov', 'www.census.gov', 'stat.gov', 'in.gov', 'www.stats.gov', 'kashi.gov', 'www.xjtj.gov', 'www.cia.gov', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.economist.com', 'books.google.com', 'www.e56.com', 'www.sbs.com', 'www.oxfordbibliographies.com', 'www.oxfordbibliographies.com', 'books.google.com', 'www.nytimes.com', 'www.reuters.com', 'books.google.com', 'www.nytimes.com', 'www.economist.com', 'thediplomat.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.google.com', 'www.technologyreview.com', 'books.google.com', 'books.google.com', 'books.google.com', 'thediplomat.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'asiatimes.com', 'books.google.com', 'world.time.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.businessinsider.com', 'www.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.theglobeandmail.com', 'books.google.com', 'books.google.com', 'indianexpress.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'apnews.com', 'www.aljazeera.com', 'books.google.com', 'books.google.com', 'www.aa.com', 'books.google.com', 'www.washingtonexaminer.com', 'books.google.com', 'books.google.com', 'www.wsj.com', 'books.google.com', 'www.businessinsider.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'china.com', 'books.google.com', 'www.todayonline.com', 'books.google.com', 'www.showcaves.com', 'www.cnn.com', 'www.google.com', 'foreignpolicy.com', 'khaleejtimes.com', 'www.latimes.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'thediplomat.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'books.google.com', 'english.peopledaily.com', 'www.wsj.com', 'www.nybooks.com', 'books.google.com', 'english.people.com', 'books.google.com', 'www.scribd.com', 'books.google.com', 'www.youtube.com', 'www.chinafile.com', 'edition.cnn.com', 'www.businessinsider.com', 'www.geopoliticalmonitor.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.google.com', 'www.courthousenews.com', 'www.businessinsider.com', 'books.google.com', 'books.google.com', 'www.reuters.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.al-monitor.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.theglobeandmail.com', 'books.google.com', 'books.google.com', 'edition.cnn.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.axios.com', 'www.youtube.com', 'foreignpolicy.com', 'www.wsj.com', 'books.google.com', 'books.google.com', 'www.google.com', 'books.google.com', 'books.google.com', 'tribune.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'news.sky.com', 'books.google.com', 'www.theartnewspaper.com', 'books.google.com', 'arabnews.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'www.britannica.com', 'www.oqya.5u.com', 'www.businessinsider.com', 'books.google.com', 'books.google.com', 'supchina.com', 'www.cnn.com', 'books.google.com', 'www.scribd.com', 'books.google.com', 'books.google.com', 'www.washingtonpost.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.meshrep.com', 'www.oed.com', 'www.nytimes.com', 'books.google.com', 'books.google.com', 'www.google.com', 'www.bbc.com', 'www.google.com', 'books.google.com', 'books.google.com', 'apnews.com', 'books.google.com', 'books.google.com', 'offbeatchina.com', 'www.voanews.com', 'www.washingtonpost.com', 'www.theartnewspaper.com', 'jamestown.org', 'www.carolinapoliticalreview.org', 'zh.wikisource.org', 'www.rfa.org', 'www.rfa.org', 'www.eastwestcenter.org', 'www.rfa.org', 'www.uyghurcongress.org', 'zh.wikisource.org', 'jamestown.org', 'www.uyghurcongress.org', 'ca.china-embassy.org', 'www.eastwestcenter.org', 'www.biblicalstudies.org', 'uyghuramerican.org', 'www.longwarjournal.org', 'newlinesinstitute.org', 'hk.plm.org', 'mesbar.org', 'hk.plm.org', 'hrw.org', 'ap.ohchr.org', 'muslimmatters.org', 'zh.wikisource.org', 'lareviewofbooks.org', 'zh.wikisource.org', 'lareviewofbooks.org', 'unesco.org', 'www.eastwestcenter.org', 'intercontinentalcry.org', ['central asian survey '], ['electrophoresis'], ['chinese journal of international law '], ['mol biol evol '], ['the journal of asian studies '], ['molecular biology and evolution'], [' inner asia ', 'brill '], ['the geographical journal'], ['americanjournal of human genetics '], ['[[bulletin of the atomic scientists'], ['refugee survey quarterly '], ['central asian survey '], ['[[rusi journal'], ['japanese journal of political science '], ['genocide studies and prevention'], ['journal of muslim minority affairs '], ['journal of medical virology '], ['journal of muslim minority affairs '], [' china quarterly '], ['genetics '], ['religion'], ['american journal of human genetics'], ['problems of post-communism '], ['scientific reports'], ['regional studies '], ['american journal of human genetics'], ['[[asian affairs'], ['journal of contemporary china '], ['open theology'], ['asian ethnicity '], ['bmc genetics'], ['bulletin of the school of oriental and african studies', 'cambridge university press on behalf of school of oriental and african studies']]",31783,Require autoconfirmed or confirmed access (no expiry set),230695,25 February 2002,Conversion script ,6203,37,2002-02-25,2002-02,2002
399,399,Campania,https://en.wikipedia.org/wiki/Campania,88,3,"['10.1093/mutage/gei076', '10.1038/nature.2016.19547', '10.2307/990664', '16434450', '26983519', None, None, None, None]","[['mutagenesis '], ['nature'], ['the journal of the society of architectural historians ']]",5,1,0,34,0,0,45,0.056818181818181816,0.011363636363636364,0.38636363636363635,0.03409090909090909,0.0,0.10227272727272728,3,"['www.av.camcom.gov', 'www.youtube.com', 'books.google.com', 'www.questia.com', 'fodors.com', 's3.amazonaws.com', 'www.thehindu.com', 'onwar.com', 'books.google.com', 'www.summerinitaly.com', 'www.oliveoilandbeyond.com', 'lifeinitaly.com', 'www.voyagesphotosmanu.com', 'www.nytimes.com', 'www.imdb.com', 'oliveoilsindia.com', 'bartleby.com', 'britannica.com', 'channel4.com', 'books.google.com', 'www.oliveoilandbeyond.com', 'www.youtube.com', 'books.google.com', 'www.youtube.com', 'www.osservatorioamianto.com', 'www.euronews.com', 'www.questia.com', 'naples.rome-in-italy.com', 'www.collinsdictionary.com', 'www.leonardocompany.com', 'naples.rome-in-italy.com', 'books.google.com', 'www.youtube.com', 'planetware.com', 'unrv.com', 'www.unesco.org', 'hdi.globaldatalab.org', 'wayback.archive-it.org', 'geonames.org', 'www.worldheritagesite.org', ['mutagenesis '], ['nature'], ['the journal of the society of architectural historians ']]",44943,Allow all users (no expiry set),80838,19 March 2002,Zisa ,1619,1,2002-03-19,2002-03,2002
400,400,Sicily,https://en.wikipedia.org/wiki/Sicily,192,4,"['10.1086/324070', '10.1515/opar-2017-0021', '10.1111/gto.12362', '10.1016/0012-821x(74)90072-7', '11573163', None, None, None, '1274378', None, None, None]","[['the american journal of human genetics '], ['open archaeology ', 'de gruyter '], ['geology today'], ['earth and planetary science letters']]",18,0,0,70,0,3,97,0.09375,0.0,0.3645833333333333,0.020833333333333332,0.0,0.11458333333333333,4,"['enel.com', 'sicilyontour.com', 'bestofsicily.com', 'historymedren.about.com', 'sicilyweb.com', 'books.google.com', 'books.google.com', 'greeknewsonline.com', 'www.initaly.com', 'porsche.com', 'britannica.com', 'books.google.com', 'italianfoodforevter.com', 'bestofsicily.com', 'britannica.com', 'books.google.com', 'books.google.com', 'fxcuisine.com', 'www.geocities.com', 'www.bestofsicily.com', 'encyclopedia.farlex.com', 'bestofsicily.com', 'www.barillaus.com', 'books.google.com', 'it.geocities.com', 'bestofsicily.com', 'bestofsicily.com', 'aboutmalta.com', 'virtuferries.com', 'www.annamariavolpi.com', 'www.bestofsicily.com', 'best-italian-wine.com', 'books.google.com', 'www.cnn.com', 'www.britannica.com', 'sicilyweb.com', 'etnavalley.com', 'thegodfathertrilogy.com', 'www.italymagazine.com', 'www.ontoeurope.com', 'knowital.com', 'books.google.com', 'bestofsicily.com', 'www.britannica.com', 'www.experiencefestival.com', 'bottlenotes.com', 'sicilyontour.com', 'bestofsicily.com', 'www.britannica.com', 'historynet.com', 'strumentires.com', 'www.ilsole24ore.com', 'books.google.com', 'www.britannica.com', 'www.italiatourismonline.com', 'books.google.com', 'books.google.com', 'www.mafia-news.com', 'www.sicilianwoodcarver.com', 'www.britannica.com', 'sicilyontour.com', 'www.wsj.com', 'www.bestofsicily.com', 'books.google.com', 'esploriamo.com', 'grifasi-sicilia.com', 'selectitaly.com', 'travelmapofsicily.com', 'grandeflanerie.com', 'italiansrus.com', 'livius.org', 'www.worldcat.org', 'storicamente.org', 'www.unesco.org', 'www.worldheritagesite.org', 'www.worldheritagesite.org', 'whc.unesco.org', 'whc.unesco.org', 'pleiades.stoa.org', 'hdi.globaldatalab.org', 'www.interamericaninstitute.org', 'www.worldheritagesite.org', 'whc.unesco.org', 'heraldica.org', 'insicilia.org', 'insicilia.org', 'whc.unesco.org', 'oah.org', ['the american journal of human genetics '], ['open archaeology ', 'de gruyter '], ['geology today'], ['earth and planetary science letters']]",27619,Require administrator access (no expiry set),156749,9 July 2001,WojPob ,6792,10,2001-07-09,2001-07,2001
401,401,Song dynasty,https://en.wikipedia.org/wiki/Song_dynasty,18,3,"['10.1038/160279b0', '10.2307/2172247', '10.1017/s0041977x13000475', None, None, None, None, None, None]","[['nature'], ['population studies'], ['bulletin of the school of oriental and african studies']]",0,0,0,3,0,0,12,0.0,0.0,0.16666666666666666,0.16666666666666666,0.0,0.16666666666666666,3,"['en.cnki.com', 'books.google.com', 'global.britannica.com', ['nature'], ['population studies'], ['bulletin of the school of oriental and african studies']]",56978,Allow all users (no expiry set),117957,9 March 2002,63.192.137.21 ,5233,6,2002-03-09,2002-03,2002
402,402,North Karnataka,https://en.wikipedia.org/wiki/North_Karnataka,33,0,[],[],3,1,0,22,0,0,7,0.09090909090909091,0.030303030303030304,0.6666666666666666,0.0,0.0,0.12121212121212122,0,"['censusindia.gov', 'www.krepublishers.com', 'www.hindu.com', 'www.hindu.com', 'articles.timesofindia.indiatimes.com', 'ourkarnataka.com', 'www.newindianexpress.com', 'www.thehindu.com', 'www.hinduonnet.com', 'www.worldstonex.com', 'www.kamat.com', 'www.craftandartisans.com', 'www.hindustantimes.com', 'www.moneycontrol.com', 'timesofindia.indiatimes.com', 'www.karnataka.com', 'ourkarnataka.com', 'www.newindianexpress.com', 'www.business-standard.com', 'www.thequint.com', 'www.kamat.com', 'www.deccanherald.com', 'www.prabhu.50g.com', 'www.metmuseum.org', 'whc.unesco.org', 'whc.unesco.org']",4685763,Allow all users (no expiry set),50184,9 April 2006,ImpuMozhi ,1595,2,2006-04-09,2006-04,2006
403,403,Sivas,https://en.wikipedia.org/wiki/Sivas,18,0,[],[],0,2,0,7,0,0,9,0.0,0.1111111111111111,0.3888888888888889,0.0,0.0,0.1111111111111111,0,"['www.mgm.gov', 'www.tcmb.gov', 'www.milliyet.com', 'books.google.com', 'books.google.com', 'www.scribd.com', 'books.google.com', 'books.google.com', 'books.google.com']",1376207,Allow all users (no expiry set),21925,9 January 2005,Llywrch ,900,0,2005-01-09,2005-01,2005
404,404,Cornish people,https://en.wikipedia.org/wiki/Cornish_people,164,6,"['10.1386/corn.19.1.60_1', '10.1386/corn.18.1.70_1', '10.1484/j.nms.3.202', None, None, None, None, None, None]","[['cornish studies ', 'university of exeter press '], ['cornish studies ', 'university of exeter press '], ['nottingham medieval studies ']]",11,13,0,8,0,0,126,0.06707317073170732,0.07926829268292683,0.04878048780487805,0.036585365853658534,0.0,0.18292682926829268,3,"['www.cornwall.gov', 'cornwall.gov', 'www.cornwall.gov', 'www.cornwall.gov', 'db.cornwall.gov', 'www.cornwall.gov', 'www.cornwall.gov', 'www.ons.gov', 'www.abs.gov', 'democracy.cornwall.gov', 'democracy.cornwall.gov', 'democracy.cornwall.gov', '2009-2017.state.gov', 'cornishstudies.com', 'www.newstatesman.com', 'artnet.com', 'krowskernewek.com', 'cornwall.com', 'www.nytimes.com', 'books.google.com', 'www.irb.com', 'www.webarchive.org', 'cornwall-opc.org', 'cornish-census2011.org', 'www.oldcornwall.org', 'www.duchyofcornwall.org', 'www.liberalhistory.org', 'www.mebyonkernow.org', 'www.flaginstitute.org', 'www.methodist-central-hall.org', 'www.mebyonkernow.org', 'www.umcwfb.org', ['cornish studies ', 'university of exeter press '], ['cornish studies ', 'university of exeter press '], ['nottingham medieval studies ']]",2300559,Allow all users (no expiry set),114328,24 July 2005,Joolz ,1869,2,2005-07-24,2005-07,2005
405,405,Ziryab,https://en.wikipedia.org/wiki/Ziryab,25,2,"['10.1163/1573-3912_islam_sim_8172', '10.1093/gmo/9781561592630.article.31002', None, None, None, None]","[['brill'], ['[[oxford university press']]",0,0,0,8,0,0,15,0.0,0.0,0.32,0.08,0.0,0.08,2,"['www.oxfordreference.com', 'books.google.com', 'archive.aramcoworld.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'almaany.com', ['brill'], ['[[oxford university press']]",2395253,Allow all users (no expiry set),20271,6 August 2005,81.178.71.128 ,907,11,2005-08-06,2005-08,2005
406,406,Malappuram district,https://en.wikipedia.org/wiki/Malappuram_district,250,3,"['10.2307/2690896', '10.1086/356288', None, None, None, None]","[['mathematics magazine '], ['isis ']]",23,50,0,112,0,0,62,0.092,0.2,0.448,0.012,0.0,0.304,2,"['censusindia.gov', 'sametham.kite.kerala.gov', 'sametham.kite.kerala.gov', 'keralapolice.gov', 'kerala.gov', 'www.censusindia.gov', 'censusindia.gov', 'spb.kerala.gov', 'www.fibkerala.gov', 'industry.kerala.gov', 'malappuram.keralapolice.gov', 'industry.kerala.gov', 'ceo.kerala.gov', 'censusindia.gov', 'delimitation.lsgkerala.gov', 'censusindia.gov', 'sametham.kite.kerala.gov', 'lsi.gov', 'homoeopathy.kerala.gov', 'censusindia.gov', 'planningcommission.gov', 'ecostat.kerala.gov', 'districts.ecourts.gov', 'sametham.kite.kerala.gov', 'lsi.gov', 'www.mlp.kerala.gov', 'lsgkerala.gov', 'ecostat.kerala.gov', 'www.ceo.kerala.gov', 'trend.kerala.gov', 'sametham.kite.kerala.gov', 'lsi.gov', 'sec.kerala.gov', 'sametham.kite.kerala.gov', 'sametham.kite.kerala.gov', 'industry.kerala.gov', 'lsgkerala.gov', 'lsgkerala.gov', 'lsgkerala.gov', 'www.ecostat.kerala.gov', 'lsi.gov', 'www.joinindiannavy.gov', 'msmedithrissur.gov', 'sametham.kite.kerala.gov', 'malappuram.keralapolice.gov', 'ecostat.kerala.gov', 'homoeopathy.kerala.gov', 'censusindia.gov', 'lsgkerala.gov', 'censusindia.gov', 'economictimes.indiatimes.com', 'www.thehindu.com', 'www.mathrubhumi.com', 'www.thehindu.com', 'books.google.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'www.deccanherald.com', 'weather.msn.com', 'www.thehindu.com', 'english.forbesmiddleeast.com', 'timesofindia.indiatimes.com', 'www.deccanchronicle.com', 'www.frontlineonnet.com', 'economictimes.indiatimes.com', 'dcbookstore.com', 'gulfnews.com', 'timesofindia.indiatimes.com', 'english.manoramaonline.com', 'www.asianage.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'epaper.malayalamvaarika.com', 'articles.timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.ethnologue.com', 'www.deccanchronicle.com', 'articles.timesofindia.indiatimes.com', 'books.google.com', 'www.mathrubhumi.com', 'www.newindianexpress.com', 'timesofindia.indiatimes.com', 'www.hindu.com', 'www.mathrubhumi.com', 'www.time.com', 'nilamburnews.com', 'www.thehindu.com', 'thenewsminute.com', 'www.onmanorama.com', 'english.mathrubhumi.com', 'www.thehindu.com', 'hellobahrain.com', 'www.hindu.com', 'rediff.com', 'www.mapsofindia.com', 'articles.timesofindia.indiatimes.com', 'www.thehindu.com', 'books.google.com', 'www.thehindu.com', 'www.mathrubhumi.com', 'www.onmanorama.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.thehindu.com', 'puzhakal0.tripod.com', 'www.ethnologue.com', 'www.thehindubusinessline.com', 'www.thehindu.com', 'post.artoflegendindia.com', 'www.deccanchronicle.com', 'www.thehindu.com', 'books.google.com', 'nativeplanet.com', 'www.thehindu.com', 'www.arabnews.com', 'www.manoramaonline.com', 'www.thehindu.com', 'touristinindia.com', 'www.hindu.com', 'nativeplanet.com', 'nwitimes.com', 'economictimes.indiatimes.com', 'www.deccanchronicle.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'nativeplanet.com', 'www.thehindu.com', 'www.vccircle.com', 'imsmagic.com', 'aryavaidyasala.com', 'nativeplanet.com', 'economictimes.indiatimes.com', 'www.ethnologue.com', 'www.newindianexpress.com', 'www.onmanorama.com', 'www.ineszupanov.com', 'articles.timesofindia.indiatimes.com', 'www.newindianexpress.com', 'www.hindu.com', 'www.variety.com', 'www.frontlineonnet.com', 'timesofindia.indiatimes.com', 'keralakaumudi.com', 'english.manoramaonline.com', 'books.google.com', 'keralartc.com', 'keralabookstore.com', 'www.nativeplanet.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.thehindu.com', 'books.google.com', 'www.hindu.com', 'www.business-standard.com', 'english.mathrubhumi.com', 'www.deccanchronicle.com', 'cnbctv18.com', 'www.keltronelcera.com', 'www.thehindu.com', 'www.financialexpress.com', 'fonts.googleapis.com', 'www.cartage.org', 'kinfra.org', 'www.malappuramtourism.org', 'keralatourism.org', 'keralasahityaakademi.org', 'keralatourism.org', 'keralatourism.org', 'naturalheritage.intach.org', 'keralatourism.org', 'keralatourism.org', 'urbanaffairskerala.org', 'malappuramtourism.org', 'keralatourism.org', 'www.keltex.org', 'malappuramtourism.org', 'en.climate-data.org', 'keralatourism.org', 'keralatourism.org', 'keralatourism.org', 'keralatourism.org', 'www.keralatourism.org', 'www.birdlife.org', 'keralatourism.org', ['mathematics magazine '], ['isis ']]",223470,Allow all users (no expiry set),241069,8 May 2003,Sudhir Krishnan~enwiki ,6063,12,2003-05-08,2003-05,2003
407,407,Palestinians,https://en.wikipedia.org/wiki/Palestinians,329,26,"['10.1086/386295', '10.1179/peq.1876.8.3.132', '10.1179/tav.1990.1990.2.223', '10.1016/j.ajhg.2017.06.013', '10.1093/molbev/msm049', '10.1111/j.1529-8817.2005.00161.x', '10.3389/fgene.2017.00087', '10.1007/s004390000426', '10.1007/s00439-003-1031-4', '10.1086/374384', '10.1371/journal.pgen.1003316', '10.1016/j.cell.2020.04.024', '10.1007/s00439-012-1235-6', '10.1179/peq.1877.9.2.89', '10.1016/j.ijintrel.2009.05.006', '10.1163/156852000511303', '10.1016/j.ajhg.2010.04.015', '10.1525/jps.1975.5.1-2.00p0373x', '10.2307/1291760', '10.1017/s0261143002002039', '10.1111/j.1354-5078.2004.00167.x', '10.3751/67.2.12', '10.1353/ncr.0.0027', '10.1016/j.fsigen.2010.08.005', '10.1038/nature09103', '10.2307/604972', '15069642', None, None, '28757201', '17351267', '15996172', '28680441', '11153918', '14586639', '12629598', '23468648', '32470400', '23052947', None, None, None, '20560205', None, None, None, None, None, None, '20843760', '20531471', None, '1181965', None, None, '5544389', None, None, '5478715', None, None, '1180338', '3585000', None, '3543766', None, None, None, '3032072', None, None, None, None, None, None, None, None, None]","[[' american journal of human genetics '], ['palestine exploration quarterly '], [' tel aviv '], ['american journal of human genetics'], [' molecular biology and evolution '], ['annals of human genetics'], ['frontiers in genetics'], ['human genetics '], ['human genetics'], ['[[american journal of human genetics'], ['plos genetics'], ['cell '], ['human genetics '], ['palestine exploration quarterly '], [' international journal of intercultural relations '], ['journal of the economic and social history of the orient '], ['[[american journal of human genetics'], ['journal of palestine studies'], ['dumbarton oaks papers'], ['popular music '], ['nations and nationalism'], ['middle east journal'], ['cr'], ['forensic science international'], ['nature'], [' journal of the american oriental society ']]",53,12,0,113,0,3,123,0.16109422492401215,0.0364741641337386,0.3434650455927052,0.0790273556231003,0.0,0.2765957446808511,26,"['www.pcbs.gov', 'www.census.gov', 'www.pcbs.gov', 'www.pcbs.gov', 'www.cbs.gov', 'mfa.gov', 'www.cbs.gov', 'www.ausstats.abs.gov', 'history.state.gov', 'www.pcbs.gov', 'www.cia.gov', 'www.pnic.gov', 'books.google.com', 'books.google.com', 'books.google.com', 'edition.cnn.com', 'books.google.com', 'museumvictoria.com', 'books.google.com', 'books.google.com', 'books.google.com', 'haaretz.com', 'thefreedictionary.com', 'books.google.com', 'books.google.com', 'www.hagar-gallery.com', 'books.google.com', 'www.britannica.com', 'www.thisweekinpalestine.com', 'books.google.com', 'www.iht.com', 'www.thisweekinpalestine.com', 'books.google.com', 'books.google.com', 'www.elsalvadorperspectives.com', 'www.iji.cgpublisher.com', 'www.maannews.com', 'www.luxner.com', 'www.saudiaramcoworld.com', 'www.al-monitor.com', 'test0.com', 'books.google.com', 'haaretz.com', 'books.google.com', 'www.ynetnews.com', 'books.google.com', 'www.ynetnews.com', 'books.google.com', 'www.thenation.com', 'books.google.com', 'www.haaretz.com', 'goliath.ecnext.com', 'books.google.com', 'books.google.com', 'www.alriyadh.com', 'www.articlearchives.com', 'food.com', 'www.reuters.com', 'api.nationalgeographic.com', 'www.themarker.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.timesofisrael.com', 'books.google.com', 'haaretz.com', 'www1.adnkronos.com', 'books.google.com', 'www.dailystar.com', 'www.foreignaffairs.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.pontas-agency.com', 'www.israelnationalnews.com', 'books.google.com', 'books.google.com', 'books.google.com', 'fortune.com', 'jewishworldreview.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'reemkelani.com', 'books.google.com', 'time.com', 'books.google.com', 'www.maannews.com', 'jpost.com', 'www.middleeastmonitor.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'jpost.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.al-monitor.com', 'books.google.com', 'www.pademographics.com', 'www.jpost.com', 'books.google.com', 'fr.jpost.com', 'www.signonsandiego.com', 'www.jordantimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.hanania.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.un.org', 'www.icj-cij.org', 'www.ps.undp.org', 'newleftreview.org', 'www.passia.org', 'www.bic.org', 'www.ameu.org', 'phonoarchive.org', 'www.meforum.org', 'domino.un.org', 'www.unhcr.org', 'www.memorialdoimigrante.org', 'www.icj-cij.org', 'www.molad.org', 'www.worldmun.org', 'www.badil.org', 'blog.palestine-studies.org', 'www.jcpa.org', 'www.encyclopedia.chicagohistory.org', 'www.nli.org', 'www.icj-cij.org', 'www.worldcat.org', 'phonoarchive.org', 'www.mideastweb.org', 'al-awdacal.org', 'www.jerusalemquarterly.org', 'domino.un.org', 'www.unrwa.org', 'www.unrwa.org', 'www.azure.org', 'www.arableagueonline.org', 'www.mideastweb.org', 'www.marxists.org', 'www.unrwa.org', 'www.pewforum.org', 'www.icj-cij.org', 'jta.org', 'www.jmcc.org', 'internal-displacement.org', 'www.un.org', 'www.al-bushra.org', 'www.azure.org', 'minorityrights.org', 'domino.un.org', 'www.unrwa.org', 'www.un.org', 'www.jmcc.org', 'odspi.org', 'repository.forcedmigration.org', 'www.erudit.org', 'www.icj-cij.org', 'www.el-funoun.org', 'www.palestinefilm.org', [' american journal of human genetics '], ['palestine exploration quarterly '], [' tel aviv '], ['american journal of human genetics'], [' molecular biology and evolution '], ['annals of human genetics'], ['frontiers in genetics'], ['human genetics '], ['human genetics'], ['[[american journal of human genetics'], ['plos genetics'], ['cell '], ['human genetics '], ['palestine exploration quarterly '], [' international journal of intercultural relations '], ['journal of the economic and social history of the orient '], ['[[american journal of human genetics'], ['journal of palestine studies'], ['dumbarton oaks papers'], ['popular music '], ['nations and nationalism'], ['middle east journal'], ['cr'], ['forensic science international'], ['nature'], [' journal of the american oriental society ']]",23267,Require administrator access (no expiry set),222324,8 October 2001,203.109.250.xxx ,8488,8,2001-10-08,2001-10,2001
408,408,Uttarandhra,https://en.wikipedia.org/wiki/Uttarandhra,29,0,[],[],0,3,0,13,0,0,13,0.0,0.10344827586206896,0.4482758620689655,0.0,0.0,0.10344827586206896,0,"['aponline.gov', 'indianculture.gov', 'core.ap.gov', 'idlebrain.com', 'www.newindianexpress.com', 'books.google.com', 'www.thehindu.com', 'www.visakhadairy.com', 'www.thehindu.com', 'www.ndtv.com', 'heavydutytravel.blogspot.com', 'www.ndtv.com', 'm.timesofindia.com', 'in.finance.yahoo.com', 'www.newindianexpress.com', 'www.ndtv.com']",10260143,Allow all users (no expiry set),31602,25 March 2007,Vgreat ,526,0,2007-03-25,2007-03,2007
409,409,Lombardy,https://en.wikipedia.org/wiki/Lombardy,104,1,"['10.1016/j.envres.2016.03.003', '26969808', None]",[['environmental research']],10,1,0,28,0,1,63,0.09615384615384616,0.009615384615384616,0.2692307692307692,0.009615384615384616,0.0,0.11538461538461539,1,"['milano.mfa.gov', 'www.cnbc.com', 'artsandculture.google.com', 'www.eupedia.com', 'www.cnn.com', 'www.iveco.com', 'www.furnishingidea.com', 'www.bbc.com', 'books.google.com', 'www.magnetimarelli.com', 'languagemonitor.com', 'www.mi-lorenteggio.com', 'www.nytimes.com', 'www.collinsdictionary.com', 'www.fondazione25aprile.com', 'www.lombardiaquotidiano.com', 'www.marketresearchreports.com', 'www.thelancet.com', 'elpais.com', 'www.gurufocus.com', 'www.iveco.com', 'www.federdoc.com', 'www.leonardocompany.com', 'www.statista.com', 'www.dutchwatersector.com', 'newsfood.com', 'www.artribune.com', 'www.mi-lorenteggio.com', 'www.leonardocompany.com', 'www-01.sil.org', 'phys.org', 'whc.unesco.org', 'whc.unesco.org', 'it.wikipedia.org', 'hdi.globaldatalab.org', 'stats.oecd.org', 'whc.unesco.org', 'whc.unesco.org', 'it.argealp.org', ['environmental research']]",43807,Allow all users (no expiry set),95181,11 March 2002,151.24.145.19 ,2200,5,2002-03-11,2002-03,2002
410,410,South East England,https://en.wikipedia.org/wiki/South_East_England,76,1,"['10.1038/217500c0', None, None]",[['nature']],8,25,0,14,0,1,27,0.10526315789473684,0.32894736842105265,0.18421052631578946,0.013157894736842105,0.0,0.4473684210526316,1,"['www.southampton.gov', 'www.medway.gov', 'www.kent.gov', 'www.dft.gov', 'www.gos.gov', 'statistics.gov', 'www.bracknell-forest.gov', 'www.education.gov', 'www.westsussex.gov', 'www.brighton-hove.gov', 'webarchive.nationalarchives.gov', 'www.rbwm.gov', 'www.ons.gov', 'www.berr.gov', 'www.statistics.gov', 'www.wokingham.gov', 'www3.hants.gov', 'www.portsmouthcc.gov', 'webarchive.nationalarchives.gov', 'www.milton-keynes.gov', 'eastsussex.gov', 'www.surreycc.gov', 'apps.oxfordshire.gov', 'www.buckscc.gov', 'www.reading.gov', 'www.uktisoutheast.com', 'www.europeantour.com', 'theconversation.com', 'docs.google.com', 'bigchurchdayout.com', 'www.icc-cricket.com', 'www.suttontrust.com', 'sciencevale.com', 'www.iwight.com', 'www.solenthotel.com', 'docs.google.com', 'www.btplc.com', 'www.newforestparishes.com', 'www.langtp.com', 'www.tnmoc.org', 'visionofbritain.org', 'www.worldcat.org', 'mas-se.org', 'www.tnmoc.org', 'wtgf.org', 'www.ashdownforest.org', 'ccskills.org', ['nature']]",52926,Allow all users (no expiry set),170365,22 May 2002,195.149.37.233 ,1138,10,2002-05-22,2002-05,2002
411,411,Culture of Montenegro,https://en.wikipedia.org/wiki/Culture_of_Montenegro,6,0,[],[],1,0,0,3,0,0,2,0.16666666666666666,0.0,0.5,0.0,0.0,0.16666666666666666,0,"['www.hollywoodreporter.com', 'mytheatrereviews.blogspot.com', 'www.britannica.com', 'www.njegos.org']",5595940,Allow all users (no expiry set),23707,16 June 2006,Conscious ,413,1,2006-06-16,2006-06,2006
412,412,Hedgehogs in culture,https://en.wikipedia.org/wiki/Hedgehogs_in_culture,8,0,[],[],1,2,0,2,0,1,2,0.125,0.25,0.25,0.0,0.0,0.375,0,"['blog.nationalarchives.gov', 'webarchive.nationalarchives.gov', 'www.fullbooks.com', 'www.mnn.com', 'www.pelister.org']",3399724,Allow all users (no expiry set),26347,12 December 2005,Cyberodin ,287,2,2005-12-12,2005-12,2005
413,413,West Africa,https://en.wikipedia.org/wiki/West_Africa,96,10,"['10.1093/acrefore/9780190277734.013.137', '10.1093/acrefore/9780190854584.013.66', '10.1146/annurev-genom-083117-021759', '10.1016/j.jasrep.2020.102658', '10.1007/bf02968406', '10.3213/1612-1651-10171', '10.1038/s41598-020-79418-4', '10.1016/j.forpol.2016.08.011', '10.1016/j.jaridenv.2016.12.011', '10.1177/2396939317739833', None, None, '29727585', None, None, None, '33431997', None, None, None, None, None, None, None, None, None, '7801626', None, None, None]","[['oxford university press'], ['oxford university press'], ['annual review of genomics and human genetics '], ['journal of archaeological science'], ['african archaeological review '], ['[[journal of african archaeology'], ['scientific reports '], ['forest policy and economics'], ['journal of arid environments '], ['international bulletin of mission research ']]",24,0,0,19,0,0,43,0.25,0.0,0.19791666666666666,0.10416666666666667,0.0,0.3541666666666667,10,"['todaygh.com', 'search.proquest.com', '--books.google.com', 'www.lonelyplanet.com', 'goal.com', 'www.nytimes.com', 'www.thoughtco.com', '--books.google.com', 'news.mongabay.com', '--books.google.com', 'www.islamreligion.com', 'www.britannica.com', 'books.google.com', 'railwaysafrica.com', 'books.google.com', 'books.google.com', 'www.bloomberg.com', 'www.lonelyplanet.com', 'books.google.com', 'www.un.org', 'www.iucn.org', 'www.imf.org', 'west-africa-brief.org', 'www.worldcat.org', 'millenniumindicators.un.org', 'nepadwatercoe.org', 'www.wipsen-africa.org', 'rainforestweb.org', 'diningforwomen.org', 'www.un.org', 'www.worldcat.org', 'www.unhcr.org', 'www.un.org', 'population.un.org', 'www.un.org', 'www.west-africa-brief.org', 'www.afdb.org', 'www.seereer.org', 'www.imf.org', 'www.uneca.org', 'unesdoc.unesco.org', 'www.mediaglobal.org', 'www.imf.org', ['oxford university press'], ['oxford university press'], ['annual review of genomics and human genetics '], ['journal of archaeological science'], ['african archaeological review '], ['[[journal of african archaeology'], ['scientific reports '], ['forest policy and economics'], ['journal of arid environments '], ['international bulletin of mission research ']]",67393,Allow all users (no expiry set),88255,3 August 2002,Jaknouse ,3063,1,2002-08-03,2002-08,2002
414,414,Brussels,https://en.wikipedia.org/wiki/Brussels,280,3,"['10.1080/09654313.2016.1139058', '10.4000/brussels.520', '10.1080/01411897908574506', None, None, None, None, None, None]","[['european planning studies', 'taylor '], ['brussels studies ', 'brussels studies [online'], ['journal of musicological research']]",14,2,0,65,0,1,195,0.05,0.007142857142857143,0.23214285714285715,0.010714285714285714,0.0,0.06785714285714285,3,"['www.state.gov', 'www.srbija.gov', 'books.google.com', 'www.euronews.com', 'books.google.com', 'www.brusselstimes.com', 'www.nytimes.com', 'www.cvent.com', 'books.google.com', 'books.google.com', 'www.stadiumguide.com', 'books.google.com', 'www.foodmuseum.com', 'books.google.com', 'books.google.com', 'www.brusselstimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'rsssf.com', 'books.google.com', 'books.google.com', 'theculturetrip.com', 'books.google.com', 'www.xpats.com', 'distcalculator.com', 'books.google.com', 'www.timesofisrael.com', 'www.nytimes.com', 'www.ft.com', 'books.google.com', 'cafébabel.com', 'books.google.com', 'books.google.com', 'www.washingtonpost.com', 'belgium.rootsweb.ancestry.com', 'books.google.com', 'books.google.com', 'city-data.com', 'eubserver.com', 'city-data.com', 'beneluxguide.com', 'books.google.com', 'www.railway-technology.com', 'www.expatistan.com', 'books.google.com', 'euobserver.com', 'books.google.com', 'guide.michelin.com', 'www.brusselstimes.com', 'euobserver.com', 'books.google.com', 'books.google.com', 'www.demographia.com', 'books.google.com', 'books.google.com', 'books.google.com', 'belgium.rootsweb.ancestry.com', 'www.fleamarketinsiders.com', 'www.brusselstimes.com', 'books.google.com', 'www.weather-atlas.com', 'books.google.com', 'www.weatherbase.com', 'uk.reuters.com', 'books.google.com', 'rsssf.com', 'www.dbnl.org', 'whc.unesco.org', 'www.dragoman.org', 'www.internations.org', 'www.foodtimeline.org', 'hdi.globaldatalab.org', 'whc.unesco.org', 'www.oecd.org', 'ich.unesco.org', 'www.vlaamsbelang.org', 'journals.openedition.org', 'whc.unesco.org', 'ich.unesco.org', 'whc.unesco.org', ['european planning studies', 'taylor '], ['brussels studies ', 'brussels studies [online'], ['journal of musicological research']]",3708,Require administrator access (no expiry set),213509,27 October 2001,203.109.250.xxx ,5813,14,2001-10-27,2001-10,2001
415,415,Montferrat,https://en.wikipedia.org/wiki/Montferrat,3,0,[],[],0,0,0,1,0,0,2,0.0,0.0,0.3333333333333333,0.0,0.0,0.0,0,['edition.cnn.com'],650849,Allow all users (no expiry set),15712,12 May 2004,Adam Bishop ,308,0,2004-05-12,2004-05,2004
416,416,Monkeys in Japanese culture,https://en.wikipedia.org/wiki/Monkeys_in_Japanese_culture,16,0,[],[],1,0,0,5,0,0,10,0.0625,0.0,0.3125,0.0,0.0,0.0625,0,"['books.google.com', 'www.sacred-texts.com', 'books.google.com', 'www.sacred-texts.com', 'books.google.com', 'openlibrary.org']",42421066,Allow all users (no expiry set),35467,6 April 2014,Keahapana ,85,2,2014-04-06,2014-04,2014
417,417,Black Forest,https://en.wikipedia.org/wiki/Black_Forest,66,0,[],[],1,0,0,9,0,0,56,0.015151515151515152,0.0,0.13636363636363635,0.0,0.0,0.015151515151515152,0,"['books.google.com', 'books.google.com', 'www.trachten-winkler.com', 'www.europeancuisines.com', 'www.britannica.com', 'pagat.com', 'www.schwarzwaldportal.com', 'www.blackforest-tourism.com', 'www.blackforeststud.com', 'www.black-forest.org']",3385,Allow all users (no expiry set),85457,24 March 2001,Rob Salzman ,1572,2,2001-03-24,2001-03,2001
418,418,Antalya,https://en.wikipedia.org/wiki/Antalya,75,1,"['10.7227/tjth.22.1.3', None, None]","[['queens college', 'the journal of transport history ']]",6,8,0,33,0,0,28,0.08,0.10666666666666667,0.44,0.013333333333333334,0.0,0.2,1,"['dergipark.gov', 'www.kgm.gov', 'dergipark.ulakbim.gov', 'www.mfa.gov', 'report.tuik.gov', 'www.mgm.gov', 'rapor.tuik.gov', 'www.antalyakulturturizm.gov', 'akmedadalya.com', 'www.kaleicimuzesi.com', 'www.likyayoluultramaratonu.com', 'hurriyetdailynews.com', 'www.milliyet.com', 'www.likyayoluultramaratonu.com', 'www.washingtontimes.com', 'secim.haberler.com', 'sabah.com', 'www.indiewire.com', 'www.sunexpress.com', 'gecce.com', 'www.ntv.com', 'kaleicimuzesi.com', 'variety.com', 'www.sabah.com', 'www.corendon-airlines.com', 'www.todayszaman.com', 'www.ucuyos.com', 'hurriyetdailynews.com', 'www.haberturk.com', 'books.google.com', 'moovitapp.com', 'independent-travellers.com', 'chpbxl.files.wordpress.com', 'www.weather2travel.com', 'moovitapp.com', 'www.weather-atlas.com', 'hurriyetdailynews.com', 'al-monitor.com', 'arama.hurriyet.com', 'sozcu.com', 'www.veooz.com', 'seatemperature.org', 'topostext.org', 'www.wdl.org', 'www.wdl.org', 'creativecommons.org', 'ant-free-zone.org', ['queens college', 'the journal of transport history ']]",361527,Allow all users (no expiry set),64158,9 November 2003,,2818,12,2003-11-09,2003-11,2003
419,419,Culture of the Basque Country,https://en.wikipedia.org/wiki/Culture_of_the_Basque_Country,3,0,[],[],0,0,0,0,0,0,3,0.0,0.0,0.0,0.0,0.0,0.0,0,[],44781105,Allow all users (no expiry set),14762,19 December 2014,Iñaki LL ,59,0,2014-12-19,2014-12,2014
420,420,İzmir,https://en.wikipedia.org/wiki/%C4%B0zmir,117,3,"['10.2307/3642952', '10.1353/hem.2004.0014', '10.2307/3643046', None, None, None, None, None, None]","[['anatolian studies ', 'british institute at ankara '], ['the hemingway review '], ['anatolian studies ', 'british institute at ankara ']]",9,8,0,45,0,0,55,0.07692307692307693,0.06837606837606838,0.38461538461538464,0.02564102564102564,0.0,0.17094017094017094,3,"['www.turkstat.gov', 'www.izmir.gov', 'www.mgm.gov', 'www.fco.gov', 'www.turkstat.gov', 'sgk.gov', 'www.sgk.gov', 'dmi.gov', 'books.google.com', 'www.webpronews.com', 'www.britannica.com', 'books.google.com', 'devlette.com', 'www.yeniasir.com', 'books.google.com', 'www.britannica.com', 'gezicini.com', 'www.adresci.com', 'books.google.com', 'www.spacecampturkey.com', 'izban.com', 'books.google.com', 'books.google.com', 'www.ds-izmir.com', 'www.eatinizmir.com', 'books.google.com', 'www.levantineheritage.com', 'gezicini.com', 'www.allaboutturkey.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.hurriyetdailynews.com', 'www.sabah.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.halkinhabercisi.com', 'kanalben.com', 'www.britannica.com', 'moovitapp.com', 'www.hastane.com', 'moovitapp.com', 'books.google.com', 'www.izban.com', 'trthaber.com', 'books.google.com', 'books.google.com', 'www.webpronews.com', 'www.ucuyos.com', 'books.google.com', 'www.aa.com', 'www.izto.org', 'www.magusa.org', 'www.akparti.org', 'dergipark.org', 'tr.m.wikipedia.org', 'climathon.climate-kic.org', 'www.npr.org', 'creativecommons.org', 'gavroche.org', ['anatolian studies ', 'british institute at ankara '], ['the hemingway review '], ['anatolian studies ', 'british institute at ankara ']]",580279,Allow all users (no expiry set),119394,6 April 2004,Llywrch ,4086,5,2004-04-06,2004-04,2004
421,421,Tourism in Algeria,https://en.wikipedia.org/wiki/Tourism_in_Algeria,41,1,"['10.1080/15583058.2015.1020458', None, None]","[['international journal of architectural heritage', '[[taylor ']]",14,2,0,13,0,0,11,0.34146341463414637,0.04878048780487805,0.3170731707317073,0.024390243902439025,0.0,0.4146341463414634,1,"['www.cia.gov', 'www.cia.gov', 'algeria.com', 'books.google.com', 'www.lemidi-dz.com', 'www.youtube.com', 'books.google.com', 'www.cliffordawright.com', 'www.algerie-focus.com', 'www.usnews.com', 'www.foodbycountry.com', 'www.lequotidien-oran.com', 'www.youtube.com', 'books.google.com', 'algeriantourism.com', 'whc.unesco.org', 'whc.unesco.org', 'whc.unesco.org', 'whc.unesco.org', 'whc.unesco.org', 'whc.unesco.org', 'www.wdl.org', 'whc.unesco.org', 'whc.unesco.org', 'whc.unesco.org', 'www.wdl.org', 'www.wdl.org', 'whc.unesco.org', 'www.discoverislamicart.org', ['international journal of architectural heritage', '[[taylor ']]",16866999,Allow all users (no expiry set),32223,10 April 2008,Anonymous101 ,271,0,2008-04-10,2008-04,2008
422,422,Minoan civilization,https://en.wikipedia.org/wiki/Minoan_civilization,201,23,"['10.1126/science.1125682', '10.1017/ccol9780521814447.014', '10.1017/s0003598x00028088', '10.1126/science.1125087', '10.1038/ncomms2871', '10.1029/2006eo340001', '10.2307/2792547', '10.1029/2006gl027205', '10.1007/bf00127003', '10.2307/630636', '10.1038/nature23310', '10.1017/s0068245400016488', '10.1017/s0003598x00079680', '10.1002/9781444355024.ch3', '10.1017/s0068245400019444', '10.9783/9781512806830-011', '10.2143/pha.20.1.3064537', '10.1007/bf00768739', '10.2972/hesp.2004.73.2.133', '10.1017/s0003581520000475', '10.1080/00438243.1998.9980386', '10.1126/science.312.5773.508', '16645092', None, None, '16645088', '23673646', None, None, None, None, None, '28783727', None, None, None, None, None, None, None, None, None, None, '16645054', None, None, None, None, '3674256', None, None, None, None, None, '5565772', None, None, None, None, None, None, None, None, None, None, None]","[['science'], ['cambridge university press'], [' antiquity '], ['science'], ['nature communications '], ['eos '], ['man '], ['geophysical research letters'], ['natural hazards'], ['the journal of hellenic studies'], ['nature'], ['the annual of the british school at athens'], [' antiquity '], ['blackwell publishing ltd '], ['the annual of the british school at athens'], ['university of pennsylvania press '], [' pharos '], ['environmental geology'], ['hesperia'], ['the antiquaries journal'], ['world archaeology '], ['science']]",17,0,0,41,0,0,120,0.0845771144278607,0.0,0.20398009950248755,0.11442786069651742,0.0,0.19900497512437812,22,"['books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.sciencedaily.com', 'books.google.com', 'www.nytimes.com', 'brewminate.com', 'books.google.com', 'wiley.com', 'books.google.com', 'university.langantiques.com', 'books.google.com', 'www.minoancrete.com', 'books.google.com', 'books.google.com', 'www.livescience.com', 'books.google.com', 'www.wired.com', 'books.google.com', 'books.google.com', 'www.fashionencyclopedia.com', 'books.google.com', 'ekathimerini.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'books.google.com', 'www.smithsonianmag.com', 'www.usatoday.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.sacred-texts.com', 'books.google.com', 'www.khanacademy.org', 'www.khanacademy.org', 'www.khanacademy.org', 'www.khanacademy.org', 'www.britishmuseum.org', 'www.agu.org', 'www.khanacademy.org', 'phys.org', 'www.therafoundation.org', 'ancient-greece.org', 'www.khanacademy.org', 'phys.org', 'www.therafoundation.org', 'arxiv.org', 'www.worldcat.org', 'www.archaeomythology.org', 'www.aegeussociety.org', ['science'], ['cambridge university press'], [' antiquity '], ['science'], ['nature communications '], ['eos '], ['man '], ['geophysical research letters'], ['natural hazards'], ['the journal of hellenic studies'], ['nature'], ['the annual of the british school at athens'], [' antiquity '], ['blackwell publishing ltd '], ['the annual of the british school at athens'], ['university of pennsylvania press '], [' pharos '], ['environmental geology'], ['hesperia'], ['the antiquaries journal'], ['world archaeology '], ['science']]",73327,Allow all users (no expiry set),120958,18 June 2002,WillWare ,4807,15,2002-06-18,2002-06,2002
423,423,Milk and meat in Jewish law,https://en.wikipedia.org/wiki/Milk_and_meat_in_Jewish_law,112,0,[],[],4,0,0,3,0,0,105,0.03571428571428571,0.0,0.026785714285714284,0.0,0.0,0.03571428571428571,0,"['books.google.com', 'www.haaretz.com', 'books.google.com', 'www.torahbase.org', 'www.sefaria.org', 'www.oqimta.org', 'www.sefaria.org']",18419834,Allow all users (no expiry set),31375,13 July 2008,Xyz7890 ,486,0,2008-07-13,2008-07,2008
424,424,Brandenburg,https://en.wikipedia.org/wiki/Brandenburg,38,1,[],[],3,0,0,4,0,1,29,0.07894736842105263,0.0,0.10526315789473684,0.02631578947368421,0.0,0.10526315789473684,0,"['en.oxforddictionaries.com', 'de.statista.com', 'de.statista.com', 'apnews.com', 'hdi.globaldatalab.org', 'commons.wikimedia.org', 'www.deutsche-metropolregionen.org']",3765,Allow all users (no expiry set),41565,1 November 2001,H. Jonat~enwiki ,1158,10,2001-11-01,2001-11,2001
425,425,Sardinia,https://en.wikipedia.org/wiki/Sardinia,219,2,"['10.1177/1464884917700914', '10.6084/m9.figshare.1263959.v5', None, None, None, None]","[['journalism'], [' figshare']]",10,1,0,29,0,0,177,0.045662100456621,0.0045662100456621,0.1324200913242009,0.0091324200913242,0.0,0.0593607305936073,2,"['weather.gov', 'www.com', 'books.google.com', 'www.cretanbeaches.com', 'www.unrv.com', 'www.kitegeneration.com', 'www.bruncuspina.com', 'www.lunarossachallenge.com', 'zanarini.wordpress.com', 'www.ilsole24ore.com', '252fwww.icis.com', 'www.news.com', 'www.avionews.com', 'earthweek.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.youtube.com', 'issuu.com', 'traveler.nationalgeographic.com', 'ethnologue.com', 'www.nonsolocinema.com', 'celtic-wrestling.tripod.com', 'www.theprimalist.com', 'www.eni.com', 'globaltwitcher.com', 'archeologianuragica.blogspot.com', 'www.rheinmetall-defence.com', 'www.aljazeera.com', 'love.sardegne.com', 'www.enricolobina.org', 'warisacrime.org', 'www.napoleon-series.org', 'www.jstor.org', 'whc.unesco.org', 'www.aristeo.org', 'pleiades.stoa.org', 'hdi.globaldatalab.org', 'eoearth.org', 'www.conifa.org', ['journalism'], [' figshare']]",29376,Allow all users (no expiry set),175517,27 December 2001,62.11.66.xxx ,4990,10,2001-12-27,2001-12,2001
426,426,"Salem, Tamil Nadu","https://en.wikipedia.org/wiki/Salem,_Tamil_Nadu",108,0,[],[],0,24,0,57,0,0,27,0.0,0.2222222222222222,0.5277777777777778,0.0,0.0,0.2222222222222222,0,"['www.salemcorporation.gov', 'www.tn.gov', 'tnpolice.gov', 'www.censusindia.gov', 'www.salemcorporation.gov', 'www.assembly.tn.gov', 'imdpune.gov', 'www.salemcorporation.gov', 'salemcorporation.gov', 'imdpune.gov', 'www.salemcorporation.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'www.tn.gov', 'cgwb.gov', 'www.indcom.tn.gov', 'www.salemcorporation.gov', 'www.assembly.tn.gov', 'www.assembly.tn.gov', 'www.salemcorporation.gov', 'www.tn.gov', 'www.assembly.tn.gov', 'archive.eci.gov', 'www.thehindu.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'collegedunia.com', 'indiamapped.com', 'www.dinakaran.com', 'www.thehindu.com', 'www.thehindu.com', 'www.tidco.com', 'www.thehindu.com', 'fallingrain.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.espncricinfo.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.thebetterindia.com', 'www.thehindu.com', 'www.thehindu.com', 'indianexpress.com', 'www.hindu.com', 'www.thehindu.com', 'www.newindianexpress.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'temple.dinamalar.com', 'www.thehindu.com', 'www.newindianexpress.com', 'www.hindu.com', 'www.thehindu.com', 'www.thehindu.com', 'www.sagoserve.com', 'www.tredyfoods.com', 'www.ndtv.com', 'www.maalaimalar.com', 'sportstar.thehindu.com', 'www.thehindu.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'airodisha.com', 'www.thehindu.com', 'www.thehindu.com', 'www.outlookindia.com', 'www.vikatan.com', 'www.thehindu.com', 'www.thehindu.com', 'www.salemmango.com', 'www.thehindu.com', 'www.thehindu.com', 'www.dnaindia.com', 'www.processregister.com', 'indianexpress.com', 'timesofindia.indiatimes.com', 'www.thehindu.com']",238919,Allow all users (no expiry set),68710,2 June 2003,Hariprasad~enwiki ,4498,0,2003-06-02,2003-06,2003
427,427,Culture of Israel,https://en.wikipedia.org/wiki/Culture_of_Israel,126,2,"['10.2307/587382', None, None]",[['the british journal of sociology']],14,6,0,61,0,0,43,0.1111111111111111,0.047619047619047616,0.48412698412698413,0.015873015873015872,0.0,0.1746031746031746,1,"['embassies.gov', 'www.galilee.gov', 'mfa.gov', 'www.mfa.gov', 'www.mfa.gov', 'www.export.gov', 'books.google.com', 'www.haaretz.com', 'www.haaretz.com', 'books.google.com', 'www.israelhayom.com', 'www.huffingtonpost.com', 'www.forward.com', 'www.israelnationalnews.com', 'www3.timeoutny.com', 'www.roberthsarkissian.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.danceinisrael.com', 'en.chessbase.com', 'books.google.com', 'en.chessbase.com', 'www.ynetnews.com', 'www.ynetnews.com', 'www.safed-kabbalah.com', 'www.britannica.com', 'www.zagraevsky.com', 'www.myjewishlearning.com', 'www.ynetnews.com', 'books.google.com', 'books.google.com', 'www.sfgate.com', 'www.highbeam.com', 'books.google.com', 'www.bloomberg.com', 'books.google.com', 'www.businessweek.com', 'www.ynetnews.com', 'www.facebook.com', 'books.google.com', 'amos-spacecom.com', 'books.google.com', 'www.lonelyplanet.com', 'books.google.com', 'nocamels.com', 'www.cbsnews.com', 'www.thejewishweek.com', 'www.nytimes.com', 'books.google.com', 'discoverymagazine.com', 'seattletimes.com', 'www.haaretz.com', 'www.myjewishlearning.com', 'www.wherefoodcomesfrom.com', 'books.google.com', 'books.google.com', 'judaism.about.com', 'books.google.com', 'ir.nasdaqomx.com', 'forward.com', 'www.travelandleisure.com', 'www.haaretz.com', 'www.britannica.com', 'www.focusmm.com', 'www.haaretz.com', 'www.hollywoodreporter.com', 'www.jewishvirtuallibrary.org', 'www.israeliconsulatela.org', 'unesdoc.unesco.org', '2fwww.olimpbase.org', 'www.jta.org', 'israel21c.org', 'www.wdl.org', 'www.parks.org', 'www.deadseascrolls.org', 'israel21c.org', 'www.jewishvirtuallibrary.org', 'www.jewishvirtuallibrary.org', 'www.jstor.org', 'www.imj.org', ['the british journal of sociology']]",211843,Allow all users (no expiry set),113901,17 April 2003,Elzamam ,1524,23,2003-04-17,2003-04,2003
428,428,Manduria,https://en.wikipedia.org/wiki/Manduria,1,0,[],[],1,0,0,0,0,0,0,1.0,0.0,0.0,0.0,0.0,1.0,0,['www.zinfandel.org'],1819879,Allow all users (no expiry set),6650,30 April 2005,Eugene van der Pijll ,108,0,2005-04-30,2005-04,2005
429,429,Tourism in San Marino,https://en.wikipedia.org/wiki/Tourism_in_San_Marino,28,1,"['10.1515/dialect-2018-0004', None, None]",[['dialectologia et geolinguistica']],4,1,0,6,0,0,16,0.14285714285714285,0.03571428571428571,0.21428571428571427,0.03571428571428571,0.0,0.21428571428571427,1,"['2009-2017.state.gov', 'www.nationalgeographic.com', 'www.visitsanmarino.com', 'www.visitsanmarino.com', 'www.inquirer.com', 'www.visitsanmarino.com', 'independent-travellers.com', 'whc.unesco.org', 'commons.wikimedia.org', 'www.worldcat.org', 'www.worldcat.org', ['dialectologia et geolinguistica']]",9023718,Allow all users (no expiry set),26366,20 January 2007,Kitia ,97,0,2007-01-20,2007-01,2007
430,430,British people,https://en.wikipedia.org/wiki/British_people,307,4,"['10.1111/j.1354-5078.1999.00053.x', '10.1093/oxfordjournals.pubjof.a029948', None, '10.1080/09662830600776694', None, None, None, None, None, None, 'govt.nz/honours/overview/honourable_privycouncil.html', None]","[['nations and nationalism'], ['publius'], [' department of the prime minister and cabinet'], ['european security']]",19,36,0,31,0,2,215,0.06188925081433225,0.11726384364820847,0.10097719869706841,0.013029315960912053,0.0,0.19218241042345277,4,"['assets.publishing.service.gov', 'scotland.gov', 'stats.gov', 'www.ons.gov', 'www.abs.gov', 'www.ons.gov', 'www.abs.gov', 'www.statssa.gov', 'nationalarchives.gov', 'factfinder.census.gov', 'abs.gov', 'nationalarchives.gov', 'www.justice.gov', 'www.statistics.gov', 'usinfo.state.gov', 'executive.gov', 'www.statssa.gov', 'www.abs.gov', 'www.royal.gov', 'www.abs.gov', 'www.london.gov', 'scotland.gov', 'www.abs.gov', 'www2.census.gov', 'www.ons.gov', 'teara.gov', 'lifeintheuktest.gov', 'state.gov', 'statistics.gov', 'itable.censtatd.gov', 'teara.gov', 'www.ons.gov', 'www.abs.gov', 'wales.gov', 'www.ons.gov', 'www.devon.gov', 'books.google.com', 'foodanddrinkeurope.com', 'books.google.com', 'statisticalatlas.com', 'encarta.msn.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'query.nytimes.com', 'tribune.com', 'books.google.com', 'www.galeon.com', 'books.google.com', 'gsy.bailiwickexpress.com', 'books.google.com', 'www.ft.com', 'sundayherald.com', 'galeon.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'worldatlas.com', 'books.google.com', 'books.google.com', 'uk.encarta.msn.com', 'hypable.com', 'books.google.com', 'theoi.com', 'uk.encarta.msn.com', 'local.live.com', 'www.itv.com', 'www.tearfund.org', 'www.ltscotland.org', 'www.thecommonwealth.org', 'electoralcommission.org', 'ippr.org', 'flaginstitute.org', 'cofe.anglican.org', 'electoralcommission.org', 'bfi.org', 'members.societe-jersiaise.org', 'assets.cambridge.org', 'catholic-ew.org', 'methodist.org', 'uup.org', 'www.solon.org', 'www.amnesty.org', 'www.mebyonkernow.org', 'visionofbritain.org', 'labour.org', ['nations and nationalism'], ['publius'], [' department of the prime minister and cabinet'], ['european security']]",19097669,Require administrator access (no expiry set),184003,21 April 2002,Fredbauder ,3930,4,2002-04-21,2002-04,2002
431,431,Negeri Sembilan,https://en.wikipedia.org/wiki/Negeri_Sembilan,46,0,[],[],0,34,0,6,0,0,6,0.0,0.7391304347826086,0.13043478260869565,0.0,0.0,0.7391304347826086,0,"['www.yns.gov', 'www.pknns.gov', 'pkwns.ns.gov', 'www.tourism.gov', 'jpsns.ns.gov', 'www.mdjl.gov', 'www.tourism.gov', 'www.mdr.gov', 'forestry.ns.gov', 'www.ns.gov', 'www.mdtampin.gov', 'muftins.gov', 'www.mppd.gov', 'www.mdkp.gov', 'www.tourism.gov', 'pmr.penerangan.gov', 'www.statistics.gov', 'nslibrary.gov', 'www.statistics.gov', 'www.mains.gov', 'www.ns.gov', 'jkrns.ns.gov', 'www.mdjl.gov', 'ptg.ns.gov', 'www.statistics.gov', 'lmns.ns.gov', 'www.mbs.gov', 'jksns.ns.gov', 'www.jkm.gov', 'jpbd.ns.gov', 'www.statistics.gov', 'pertanian.ns.gov', 'dvsns.ns.gov', 'jheains.ns.gov', 'go2travelmalaysia.com', 'www.nilaimc.com', 'books.google.com', 'www.columbiaasia.com', 'museumvolunteersjmm.com', 'www.ssh.kpjhealth.com']",376437,Allow all users (no expiry set),38243,23 November 2003,Jpatokal ,820,2,2003-11-23,2003-11,2003
432,432,Macedonia (ancient kingdom),https://en.wikipedia.org/wiki/Macedonia_(ancient_kingdom),492,4,"['10.1086/671786', '10.2307/630417', '10.4467/20834624sl.16.006.5152', '10.2307/1170959', None, None, None, None, None, None, None, None]","[[' classical philology ', 'the [[university of chicago press'], ['the journal of hellenic studies'], ['studia linguistica universitatis iagellonicae cracoviensis '], ['social science history']]",2,0,0,61,0,0,425,0.0040650406504065045,0.0,0.12398373983739837,0.008130081300813009,0.0,0.012195121951219513,4,"['books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.seeker.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'sino-platonic.org', 'www.livius.org', [' classical philology ', 'the [[university of chicago press'], ['the journal of hellenic studies'], ['studia linguistica universitatis iagellonicae cracoviensis '], ['social science history']]",42012,Require administrator access (no expiry set),221909,26 February 2002,David Parker ,4010,1,2002-02-26,2002-02,2002
433,433,Novi Sad,https://en.wikipedia.org/wiki/Novi_Sad,80,0,[],[],6,11,0,16,0,0,47,0.075,0.1375,0.2,0.0,0.0,0.2125,0,"['stat.gov', 'www.mp.gov', 'stat.gov', 'webrzs.stat.gov', 'www.puma.vojvodina.gov', 'stat.gov', 'www.hidmet.gov', 'www.hidmet.gov', 'stat.gov', 'pod2.stat.gov', 'stat.gov', 'www.bbc.com', 'www.irishnews.com', 'books.google.com', 'kanal9ns.com', 'www.coolhunting.com', 'www.nsfair.com', 'ekapija.com', 'books.google.com', 'www.eurofencingns2018.com', 'theculturetrip.com', 'www.hungarianquarterly.com', 'www.bbc.com', 'www.linguasport.com', 'www.rpkns.com', 'www.nacionalnarevija.com', 'www.mojnovisad.com', 'climate-data.org', 'meteo-climat-bzh.dyndns.org', 'www.dkv.org', 'www.novisadtourism.org', 'eng.exitfest.org', 'www.psdzeleznicarns.org']",113288,Allow all users (no expiry set),85754,19 October 2002,18.252.2.32 ,4058,11,2002-10-19,2002-10,2002
434,434,Bengali Muslims,https://en.wikipedia.org/wiki/Bengali_Muslims,159,3,"['10.1080/00856400802192952', '10.1080/14608940801997218', '10.1177/097194580400700101', None, None, None, None, None, None]","[[' south asia'], ['national identities '], [' the medieval history journal']]",36,5,0,67,0,0,48,0.22641509433962265,0.031446540880503145,0.42138364779874216,0.018867924528301886,0.0,0.27672955974842767,3,"['dl.nlb.gov', 'www.ons.gov', '2009-2017.state.gov', 'www.censusindia.gov', 'www.railway.gov', 'www.aljazeera.com', 'www.aljazeera.com', 'books.google.com', 'www.cambridgescholars.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'indianexpress.com', 'www.dhakatribune.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'worldpopulationreview.com', 'm.economictimes.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'global.britannica.com', 'www.washingtontimes.com', 'archive.dhakatribune.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.hindustantimes.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'indianexpress.com', 'filmfare.com', 'usatoday30.usatoday.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.bangladesh-web.com', 'www.hindustantimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'bqdoha.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'abc-clio.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'news.webindia123.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.bbc.com', 'books.google.com', 'en.banglapedia.org', 'en.banglapedia.org', 'en.banglapedia.org', 'en.banglapedia.org', 'www.iranicaonline.org', 'en.banglapedia.org', 'en.banglapedia.org', 'en.banglapedia.org', 'nobelprize.org', 'en.banglapedia.org', 'irfi.org', 'en.banglapedia.org', 'en.banglapedia.org', 'www.bmri.org', 'en.banglapedia.org', 'en.banglapedia.org', 'alalodulal.org', 'pewforum.org', 'alalodulal.org', 'en.banglapedia.org', 'iranicaonline.org', 'en.banglapedia.org', 'en.banglapedia.org', 'publishing.cdlib.org', 'en.banglapedia.org', 'bea-bd.org', 'www.globalreligiousfutures.org', 'en.banglapedia.org', 'en.banglapedia.org', 'en.banglapedia.org', 'en.banglapedia.org', 'en.banglapedia.org', 'www.migrationpolicy.org', 'en.banglapedia.org', 'publishing.cdlib.org', 'www.un.org', [' south asia'], ['national identities '], [' the medieval history journal']]",41787383,Allow all users (no expiry set),92384,30 January 2014,Messiaindarain ,1158,15,2014-01-30,2014-01,2014
435,435,Icelanders,https://en.wikipedia.org/wiki/Icelanders,73,16,"['10.1086/302816', '10.1126/science.aar2625', '10.2307/3005071', '10.1111/1467-8322.00023', '10.1126/science.306.5700.1278', '10.1136/bmj.319.7207.441', '10.1515/njmr-2017-0012', '10.2307/2173366', '10.1111/j.1468-0289.1957.tb00672.x', '10.1038/78036', '10.2307/3004589', '10.1086/303046', '10.2307/2886763', '10.1111/j.1467-8306.1963.tb00454.x', '10.1038/s41588-017-0031-6', '10.1002/ajpa.21419', '10712214', '29853688', None, None, '15550636', '10445931', None, '11630504', None, '10932173', None, '10931763', None, None, '29335549', '21069749', '1288180', None, None, None, None, '1127047', None, None, None, None, None, '1287529', None, None, None, None]","[[' american journal of human genetics '], ['science '], ['journal of social forces '], ['anthropology today '], ['science '], [' bmj '], [' nordic journal of migration research '], ['population studies '], ['the economic history review '], ['nature genetics '], ['social forces '], ['am. j. hum. genet. '], ['speculum '], ['annals of the association of american geographers '], [' nature genetics '], ['am. j. phys. anthropol. ']]",3,3,0,8,0,0,43,0.0410958904109589,0.0410958904109589,0.1095890410958904,0.2191780821917808,0.0,0.3013698630136986,16,"['memory.loc.gov', 'dfat.gov', 'factfinder.census.gov', 'www.electricscotland.com', 'books.google.com', 'books.google.com', 'irishtimes.com', 'www.washingtonisland.com', 'www.usaweekend.com', 'books.google.com', 'www.nationalgeographic.com', 'www.genomenewsnetwork.org', 'www.faqs.org', 'www.un.org', [' american journal of human genetics '], ['science '], ['journal of social forces '], ['anthropology today '], ['science '], [' bmj '], [' nordic journal of migration research '], ['population studies '], ['the economic history review '], ['nature genetics '], ['social forces '], ['am. j. hum. genet. '], ['speculum '], ['annals of the association of american geographers '], [' nature genetics '], ['am. j. phys. anthropol. ']]",832158,Require administrator access (no expiry set),43077,16 July 2004,Saforrest ,996,3,2004-07-16,2004-07,2004
436,436,Arroz a la valenciana,https://en.wikipedia.org/wiki/Arroz_a_la_valenciana,18,0,"[None, None, None]","[['revista d', 'departament de cultura de la generalitat de catalunya']]",1,0,0,11,0,0,5,0.05555555555555555,0.0,0.6111111111111112,0.0,0.0,0.05555555555555555,1,"['www.degustalarioja.com', 'books.google.com', 'epoca1.valenciaplaza.com', 'books.google.com', 'cadenaser.com', 'gastronomiabolivia.com', 'recetasdenicaragua.com', 'elcomidista.elpais.com', 'www.elmundotoday.com', 'hispanoplaces.com', 'www.geocities.com', 'www.worldcat.org', ['revista d', 'departament de cultura de la generalitat de catalunya']]",10226955,Allow all users (no expiry set),15460,23 March 2007,LaNicoya ,132,1,2007-03-23,2007-03,2007
437,437,Ponnani,https://en.wikipedia.org/wiki/Ponnani,54,0,[],[],4,11,0,9,0,0,30,0.07407407407407407,0.2037037037037037,0.16666666666666666,0.0,0.0,0.2777777777777778,0,"['censusindia.gov', 'censusindia.gov', 'lsi.gov', 'www.ponnanimunicipality.lsgkerala.gov', 'sec.kerala.gov', 'lsgkerala.gov', 'malappuram.keralapolice.gov', 'lsgkerala.gov', 'censusindia.gov', 'malappuram.keralapolice.gov', 'dgllnoida.gov', 'www.thehindu.com', 'travel.manoramaonline.com', 'www.mathrubhumi.com', 'books.google.com', 'www.arabnews.com', 'www.hindu.com', 'www.hindu.com', 'www.ineszupanov.com', 'nativeplanet.com', 'www.cartage.org', 'malappuramtourism.org', 'www.keralatourism.org', 'www.mesponnanicollege.org']",3087764,Allow all users (no expiry set),49911,5 November 2005,SHYAM b1281 ,761,2,2005-11-05,2005-11,2005
438,438,Tamil Muslim,https://en.wikipedia.org/wiki/Tamil_Muslim,32,2,"['10.1093/jis/2.1.25', 'abs/10.1080/13602009708716375?journalcode=cjmm20', '15455059', None, '355923', None]","[['journal of islamic studies'], ['journal of muslim minority affairs', '[[journal of muslim minority affairs']]",1,0,0,14,0,0,15,0.03125,0.0,0.4375,0.0625,0.0,0.09375,2,"['hindu.com', 'www.india.com', 'books.google.com', 'littleindia.com', 'books.google.com', 'www.thehindu.com', 'hindu.com', 'www.hanafionline.com', 'frontline.thehindu.com', 'books.google.com', 'www.hindu.com', 'www.islamicvoice.com', 'ier.sagepub.com', 'www.thehindu.com', 'www.countercurrents.org', ['journal of islamic studies'], ['journal of muslim minority affairs', '[[journal of muslim minority affairs']]",3095462,Allow all users (no expiry set),20206,6 November 2005,202.56.231.116 ,1808,10,2005-11-06,2005-11,2005
439,439,Yorkshire,https://en.wikipedia.org/wiki/Yorkshire,279,1,[],[],36,11,0,67,0,9,156,0.12903225806451613,0.03942652329749104,0.24014336917562723,0.0035842293906810036,0.0,0.17204301075268819,0,"['www.countryside.gov', 'www.statistics.gov', 'www.statistics.gov', 'www.york.gov', 'www.legislation.gov', 'www.kirklees.gov', 'www.countryside.gov', 'www.wakefield.gov', 'www.york.gov', 'www.highways.gov', 'www.opsi.gov', 'sheffieldfc.com', 'moovitapp.com', 'www.shadowdrake.com', 'fortunecity.com', 'northernlifestyle.com', 'www.britaingallery.com', 'books.google.com', 'www.studyyorkshire.com', 'www.theknowledgeonline.com', 'moovitapp.com', 'www.fifa.com', 'www.yorkshire.com', 'conservatives.com', 'www.youtube.com', 'fileybay.com', 'britannia.com', 'www.historic-uk.com', 'books.google.com', 'everything.com', 'aboutfood.com', 'crwflags.com', 'britainexpress.com', 'www.fifa.com', 'dracula-in-whitby.com', 'boozecruise.com', 'www.simonarmitage.com', 'books.google.com', 'www.bbc.com', 'britainexpress.com', 'britainexpress.com', 'w.fixtureslive.com', 'artchive.com', 'www.etymonline.com', 'robinhoodairport.com', 'www.premiershiprugby.com', 'history-timeline.deepthi.com', 'www.yorkshire-forward.com', 'britannia.com', 'about.com', 'www.uefa.com', 'yorkshirehistory.com', 'ifhof.com', 'beer-pages.com', 'digyorkshire.com', 'books.google.com', 'www.britainexpress.com', 'airports-worldwide.com', 'www.imdb.com', 'summer-wine.com', 'www.time.com', 'digyorkshire.com', 'news.sky.com', 'www.britainexpress.com', 'www.radiotimes.com', 'in.news.yahoo.com', 'worlds.yorkshire.com', 'books.google.com', 'seymour-recipes.com', 'www.visitbradford.com', 'www.youtube.com', 'books.google.com', 'books.google.com', 'www.rugbypass.com', 'knotfest.com', 'www.nytimes.com', 'www.yorkromanfestival.com', 'richardiii.com', 'creativecommons.org', 'www.yorkshireha.org', 'num.org', 'www.naturalengland.org', 'brontefamily.org', 'www.arch.wyjs.org', 'www.conifa.org', 'newadvent.org', 'oneyorkshire.org', 'thoresby.org', 'www.churchofengland.org', 'www.yorkshiredialectsociety.org', 'universalteacher.org', 'wensleydale.org', 'sqa.org', 'genuki.org', 'theotherpages.org', 'www.nationaltrust.org', 'www.visityork.org', 'localhistories.org', 'www.iht.org', 'romans-in-britain.org', 'www.english-heritage.org', 'yorkshireawards.org', 'www.visionofbritain.org', 'haworth-village.org', 'rspb.org', 'genuki.org', 'rlhalloffame.org', 'www.yorkshireridings.org', 'lgbce.org', 'quaffale.org', 'visityork.org', 'rlhalloffame.org', 'nrm.org', 'luminarium.org']",36637,Allow all users (no expiry set),192216,26 January 2002,MichaelTinkler ,4046,6,2002-01-26,2002-01,2002
440,440,Alsace,https://en.wikipedia.org/wiki/Alsace,35,0,[],[],2,0,0,6,0,0,27,0.05714285714285714,0.0,0.17142857142857143,0.0,0.0,0.05714285714285714,0,"['books.google.com', 'books.google.com', 'global.oup.com', 'timesmachine.nytimes.com', 'bellefrance.com', 'books.google.com', 'www.britishcouncil.org', 'www.unserland.org']",48129,Allow all users (no expiry set),84375,7 April 2002,Pgdudda ,2800,10,2002-04-07,2002-04,2002
441,441,Wallonia,https://en.wikipedia.org/wiki/Wallonia,68,1,"['10.3406/rnord.1962.2410', None, None]",[['revue du nord']],0,2,0,12,0,0,53,0.0,0.029411764705882353,0.17647058823529413,0.014705882352941176,0.0,0.04411764705882353,1,"['www.cia.gov', 'sos.maryland.gov', 'www.answers.com', 'books.google.com', 'artsandfaith.com', 'artnet.com', 'www.world-gazetteer.com', 'books.google.com', 'allstates-flag.com', 'efi-costarica.com', 'practicallyedible.com', 'theage.com', 'etymonline.com', 'etymonline.com', ['revue du nord']]",99721,Allow all users (no expiry set),72294,5 October 2002,Montrealais ,2484,4,2002-10-05,2002-10,2002
442,442,Culture of Kathmandu,https://en.wikipedia.org/wiki/Culture_of_Kathmandu,14,0,[],[],2,3,0,3,0,0,6,0.14285714285714285,0.21428571428571427,0.21428571428571427,0.0,0.0,0.35714285714285715,0,"['www.kathmandu.gov', 'www.kathmandu.gov', 'nepal.usembassy.gov', 'www.asiatravel.com', 'www.asiatravel.com', 'www.nepalitimes.com', 'www.aarohantheatre.org', 'kathmanduarts.org']",32227770,Allow all users (no expiry set),27481,27 June 2011,Dr. Blofeld ,72,0,2011-06-27,2011-06,2011
443,443,Sabah,https://en.wikipedia.org/wiki/Sabah,552,13,"['10.2307/851525', '10.1017/s0022463401000042', '10.1579/05-s-093.1', '10.4000/moussons.3454', '10.4249/scholarpedia.1', '10.2307/2642463', '10.1111/j.1365-2699.2009.02243.x', '10.1108/jmd-02-2015-0019', '10.1029/2007jd009218', '10.3406/arch.1999.3538', '10.1177/0967828x9600400105', '10.1353/cch.2007.0009', '10.1155/2013/358183', None, None, '16989512', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None]","[[' ethnomusicology'], ['journal of southeast asian studies '], ['ambio '], [' social science research on southeast asia'], ['scholarpedia ', 'public works department '], [' asian survey'], ['institute for tropical biology and conservation'], ['universiti teknologi mara'], [' journal of geophysical research'], ['archipel '], [' south east asia research'], ['journal of colonialism and colonial history '], ['journal of ecosystems ']]",38,74,0,367,0,2,62,0.06884057971014493,0.13405797101449277,0.6648550724637681,0.02355072463768116,0.0,0.22644927536231885,13,"['www.ww2australia.gov', 'www.dmpm.nre.gov', 'dfa.gov', 'eresources.nlb.gov', 'www.sabah.gov', 'www.dosm.gov', 'www.ssl.sabah.gov', 'discovery.nationalarchives.gov', 'www.kpi.sabah.gov', 'dfa.gov', 'www.mot.gov', 'ww2.sabah.gov', 'jpnsabah.moe.gov', 'ww2.sabah.gov', 'tvi.rtm.gov', 'www.pusat-sejarah.gov', 'www.skmm.gov', 'ww2.sabah.gov', 'www.dosm.gov', 'www.dvs.gov', 'ww2.sabah.gov', 'sabahvfm.rtm.gov', 'discovery.nationalarchives.gov', 'sabahfm.rtm.gov', 'www.forest.sabah.gov', 'museum.sabah.gov', 'www.wildlife.sabah.gov', 'www.legislation.gov', 'rmk11.epu.gov', 'www.sabah.gov', 'www.statistics.gov', 'eresources.nlb.gov', 'www.awm.gov', 'www.awm.gov', 'www.did.sabah.gov', 'www.idfr.gov', 'www.museum.sabah.gov', 'emisportal.moe.gov', 'www.lawnet.sabah.gov', 'etp.pemandu.gov', 'rmk11.epu.gov', 'www.deped.gov', 'www.officialgazette.gov', 'www.dosm.gov', 'pmr.penerangan.gov', 'corporate.tourism.gov', 'www.sabah.gov', 'www.lawnet.sabah.gov', 'ww2.sabah.gov', 'mvc.gov', 'www.jpn.gov', 'www.sabah.gov', 'www.msn.sabah.gov', 'eresources.nlb.gov', 'ww2.sabah.gov', 'www.sabah.gov', 'etp.pemandu.gov', 'www.sabah.gov', 'lpps.sabah.gov', 'www.fishdept.sabah.gov', 'www.lawnet.sabah.gov', 'www.lawnet.sabah.gov', 'www.dosm.gov', 'www.mot.gov', 'www.bbec.sabah.gov', 'www.awm.gov', 'www.statistics.gov', 'www.sabah.gov', 'www.sabah.gov', 'ww2.sabah.gov', 'www.statistics.gov', 'trove.nla.gov', 'www.lpps.sabah.gov', 'ww2.sabah.gov', 'books.google.com', 'www.theborneopost.com', 'books.google.com', 'www.sinarharian.com', 'www.freemalaysiatoday.com', 'www.malaysianwireless.com', 'books.google.com', 'kk12fm.com', 'www.thestar.com', 'www.nestle.com', 'news.abs-cbn.com', 'www.theborneopost.com', 'www.thestar.com', 'www.theborneopost.com', 'articles.chicagotribune.com', 'books.google.com', 'books.google.com', 'www.etawau.com', 'books.google.com', 'www.straitstimes.com', 'www.theborneopost.com', 'www.newsarawaktribune.com', 'books.google.com', 'farm8.staticflickr.com', 'news.google.com', 'www.theborneopost.com', 'books.google.com', 'books.google.com', 'marimariculturalvillage.com', 'www.theborneopost.com', 'malaysiandigest.com', 'www.theborneopost.com', 'www.questia.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.economist.com', 'www.etawau.com', 'books.google.com', 'www.dailyexpress.com', 'books.google.com', 'www.philstar.com', 'www.theborneopost.com', 'says.com', 'www.highbeam.com', 'borneobulletin.com', 'books.google.com', 'www.thestar.com', 'books.google.com', 'www.freemalaysiatoday.com', 'www.antarasulteng.com', 'www.utusan.com', 'www.themalaymailonline.com', 'books.google.com', 'dailyexpress.com', 'm.themalaymailonline.com', 'www.thestar.com', 'books.google.com', 'www.mindanews.com', 'books.google.com', 'www.dailyexpress.com', 'www.theborneopost.com', 'www.dailyexpress.com', 'www.thestar.com', 'www.theborneopost.com', 'www.bharian.com', 'books.google.com', 'books.google.com', 'www.thestar.com', 'www.dailyexpress.com', 'www.etawau.com', 'www.theborneopost.com', 'www.thestar.com', 'books.google.com', 'books.google.com', 'www.newsabahtimes.com', 'www.nst.com', 'books.google.com', 'www.dailyexpress.com', 'www.thestar.com', 'www.dailyexpress.com', 'books.google.com', 'www.dailyexpress.com', 'www.dailyexpress.com', 'www.themalaymailonline.com', 'says.com', 'books.google.com', 'books.google.com', 'www.therakyatpost.com', 'www.theborneopost.com', 'www.astroawani.com', 'books.google.com', 'www.pressreader.com', 'books.google.com', 'www.borneolegend.com', 'www.theglobeandmail.com', 'news.google.com', 'news.google.com', 'www.kkfoodfest.com', 'books.google.com', 'www.dailyexpress.com', 'www.nst.com', 'books.google.com', 'books.google.com', 'www.thestar.com', 'www.dailyexpress.com', 'www.dailyexpress.com', 'www.dailyexpress.com', 'kkjazzfest.com', 'www.thestar.com', 'youtube.com', 'www.theborneopost.com', 'books.google.com', 'books.google.com', 'www.theborneopost.com', 'books.google.com', 'ww1.utusan.com', 'youtube.com', 'www.thestar.com', 'www.themalaymailonline.com', 'cybo.com', 'www.sunstar.com', 'www.thestar.com', 'dailyexpress.com', 'books.google.com', 'www.sabahfest.com', 'news.google.com', 'www.rsssf.com', 'books.google.com', 'www.newsabahtimes.com', 'books.google.com', 'books.google.com', 'www.thestar.com', 'books.google.com', 'books.google.com', 'www.sedia.com', 'news.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.dailyexpress.com', 'www.dailyexpress.com', 'www.theborneopost.com', 'www.straitstimes.com', 'www.nst.com', 'www.bernama.com', 'www.nst.com', 'www.theborneopost.com', 'www.nst.com', 'www.straitstimes.com', 'm.themalaymailonline.com', 'www.dailyexpress.com', 'travel.asiaone.com', 'www.theborneopost.com', 'www.skyscanner.com', 'www.theborneopost.com', 'cybo.com', 'books.google.com', 'news.google.com', 'www.thestar.com', 'malaysiandigest.com', 'doesitsnowin.com', 'www.sinchew.com', 'www.therakyatpost.com', 'books.google.com', 'www.dailyexpress.com', 'books.google.com', 'www.thejakartapost.com', 'www.theborneopost.com', 'dailyexpress.com', 'www.thestar.com', 'books.google.com', 'books.google.com', 'www.dailyexpress.com', 'dailyexpress.com', 'books.google.com', 'www.malaymail.com', 'books.google.com', 'www.seatrade-maritime.com', 'books.google.com', 'books.google.com', 'books.google.com', 'traveltips.usatoday.com', 'cybo.com', 'books.google.com', 'palawan-news.com', 'www.dailyexpress.com', 'www.suriagroup.com', 'www.vokfmsabah.com', 'www.nst.com', 'www.theborneopost.com', 'books.google.com', 'books.google.com', 'www.dailyexpress.com', 'm.detik.com', 'www.theborneopost.com', 'www.newsabahtimes.com', 'www.dailyexpress.com', 'jesseltonpoint.com', 'books.google.com', 'www.dailyexpress.com', 'www.thestar.com', 'books.google.com', 'www.thestar.com', 'www.therakyatpost.com', 'www.freemalaysiatoday.com', 'www.malaymail.com', 'www.nytimes.com', 'www.irishtimes.com', 'www.dailyexpress.com', 'www.dailyexpress.com', 'www.themalaymailonline.com', 'www.theborneopost.com', 'www.dailyexpress.com', 'books.google.com', 'www.dailyexpress.com', 'www.geoexpro.com', 'www.dailyexpress.com', 'books.google.com', 'www.dailyexpress.com', 'www.bworldonline.com', 'www.newsabahtimes.com', 'www.dailyexpress.com', 'www.theborneopost.com', 'books.google.com', 'books.google.com', 'dailyexpress.com', 'themalaysianreserve.com', 'books.google.com', 'books.google.com', 'www.theborneopost.com', 'news.google.com', 'www.thestar.com', 'www.dailyexpress.com', 'www.theborneopost.com', 'www.oxfordbusinessgroup.com', 'www.sabahnewstoday.com', 'books.google.com', 'www.theborneopost.com', 'www.dailyexpress.com', 'www.themalaymailonline.com', 'books.google.com', 'www.theborneopost.com', 'www.dailyexpress.com', 'books.google.com', 'www.malaysiandigest.com', 'www.dailyexpress.com', 'www.gmanetwork.com', 'www.dailyexpress.com', 'www.therakyatpost.com', 'books.google.com', 'www.theborneopost.com', 'www.theborneopost.com', 'dailyexpress.com', 'books.google.com', 'www.theborneopost.com', 'www.dailyexpress.com', 'books.google.com', 'www.reuters.com', 'www.dailyexpress.com', 'www.theborneopost.com', 'www.thestar.com', 'www.dailyexpress.com', 'safarimuseum.com', 'www.grin.com', 'www.theborneopost.com', 'books.google.com', 'www.newsabahtimes.com', 'www.flyingdusun.com', 'news.google.com', 'www.sabahtourism.com', 'www.mb.com', 'news.google.com', 'borneobulletin.com', 'books.google.com', 'www.thestar.com', 'books.google.com', 'news.google.com', 'www.businesscircle.com', 'www.theantdaily.com', 'www.thestar.com', 'books.google.com', 'says.com', 'news.mb.com', 'books.google.com', 'books.google.com', 'news.google.com', 'www.malaysiandigest.com', 'books.google.com', 'www.etawau.com', 'books.google.com', 'books.google.com', 'tv.com', 'www.soyacincau.com', 'books.google.com', 'books.google.com', 'www.theborneopost.com', 'books.google.com', 'www.thestar.com', 'books.google.com', 'www.thestar.com', 'www.highbeam.com', 'www.theedgemarkets.com', 'news.google.com', 'www.ocdn.com', 'www.dailyexpress.com', 'books.google.com', 'www.bt.com', 'books.google.com', 'books.google.com', 'www.thestar.com', 'www.theborneopost.com', 'borneobulletin.com', 'books.google.com', 'news.google.com', 'news.mongabay.com', 'www.theborneopost.com', 'www.dailyexpress.com', 'www.malaymail.com', 'www.thestar.com', 'www.theborneopost.com', 'www.dailyexpress.com', 'www.sabahair.com', 'books.google.com', 'www.themalaymailonline.com', 'www.bt.com', 'www.borneobirdfestival.com', 'www.bt.com', 'www.dailyexpress.com', 'www.astroawani.com', 'upsidedownhouse.com', 'www.bt.com', 'www.dailyexpress.com', 'www.oxfordbusinessgroup.com', 'www.e-borneo.com', 'books.google.com', 'books.google.com', 'www.malaysiandigest.com', 'www.bbc.com', 'www.theborneopost.com', 'books.google.com', 'www.flyingdusun.com', 'www.asiaone.com', 'www.newsabahtimes.com', 'www.newsabahtimes.com', 'www.sedia.com', 'www.dailyexpress.com', 'books.google.com', 'www.astro.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.channelnewsasia.com', 'books.google.com', 'www.suteraharbour.com', 'news.google.com', 'books.google.com', 'www.thestar.com', 'books.google.com', 'www.thestar.com', 'm.themalaymailonline.com', 'sea.mashable.com', 'www.newsabahtimes.com', 'www.upsidedownhouse.com', 'news.google.com', 'www.pressreader.com', 'wwf.panda.org', 'www.gutenberg.org', 'www.ccel.org', 'www.commonlii.org', 'foreversabah.org', 'www.bsbcc.org', 'www.newmandala.org', 'www.ocasia.org', 'treaties.un.org', 'www.ijssh.org', 'www.bsbcc.org', 'www.seaa-web.org', 'www.un.org', 'rsis.ramsar.org', 'www.sabahparks.org', 'www.icj-cij.org', 'amti.csis.org', 'hdi.globaldatalab.org', 'www.yayasansabahgroup.org', 'planipolis.iiep.unesco.org', 'wwf.panda.org', 'treaties.un.org', 'www.fao.org', 'www.csis.org', 'www.my.undp.org', 'www.sabahparks.org', 'www.sino-platonic.org', 'asiafoundation.org', 'www.sabahparks.org', 'treaties.un.org', 'www.unodc.org', 'www.newmandala.org', 'www.beff.org', 'www.sabahparks.org', 'whc.unesco.org', 'www.un.org', 'foreversabah.org', 'www.gsm.org', [' ethnomusicology'], ['journal of southeast asian studies '], ['ambio '], [' social science research on southeast asia'], ['scholarpedia ', 'public works department '], [' asian survey'], ['institute for tropical biology and conservation'], ['universiti teknologi mara'], [' journal of geophysical research'], ['archipel '], [' south east asia research'], ['journal of colonialism and colonial history '], ['journal of ecosystems ']]",28678,Allow all users (no expiry set),334902,28 October 2001,195.149.37.xxx ,5364,6,2001-10-28,2001-10,2001
444,444,Beary,https://en.wikipedia.org/wiki/Beary,49,0,[],[],1,4,0,28,0,0,16,0.02040816326530612,0.08163265306122448,0.5714285714285714,0.0,0.0,0.10204081632653061,0,"['catalog.loc.gov', 'catalog.loc.gov', 'catalog.loc.gov', 'catalog.loc.gov', 'www.daijiworld.com', 'www.flickr.com', 'www.daijiworld.com', 'www.deccanherald.com', 'hindu.com', 'www.coastaldigest.com', 'www.daijiworld.com', 'hindu.com', 'www.daijiworld.com', 'www.daijiworld.com', 'mangalorean.com', 'www.thehindu.com', 'www.daijiworld.com', 'www.daijiworld.com', 'www.daijiworld.com', 'www.ksajonline.com', 'www.daijiworld.com', 'www.coastaldigest.com', 'www.daijiworld.com', 'www.daijiworld.com', 'www.mangaloretoday.com', 'www.coastaldigest.com', 'www.daijiworld.com', 'www.thenewsminute.com', 'www.daijiworld.com', 'www.daijiworld.com', 'www.daijiworld.com', 'www.kannadigaworld.com', 'www.salafiksa.org']",4683805,Allow all users (no expiry set),36869,9 April 2006,Lordshaneez ,1341,1,2006-04-09,2006-04,2006
445,445,Coimbatore,https://en.wikipedia.org/wiki/Coimbatore,310,1,"['10.11609/jott.zpj.1657.2944-8', None, None]",[['zoos']],7,33,0,218,0,0,51,0.02258064516129032,0.1064516129032258,0.7032258064516129,0.0032258064516129032,0.0,0.13225806451612904,1,"['imdpune.gov', 'www.tn.gov', 'www.censusindia.gov', 'archive.eci.gov', 'imdpune.gov', 'www.censusindia.gov', 'www.tn.gov', 'censusindia.gov', 'www.tn.gov', 'eservices.tnpolice.gov', 'pibmumbai.gov', 'www.censusindia.gov', 'payment.ccmc.gov', 'censusindia.gov', 'www.censusindia.gov', 'censusindia.gov', 'allindiaradio.gov', 'ifgtb.icfre.gov', 'www.ccmc.gov', 'censusindia.gov', 'www.censusindia.gov', 'allindiaradio.gov', 'pib.gov', 'censusindia.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'www.ncrb.gov', 'moud.gov', 'www.indianrail.gov', 'www.ccmc.gov', 'www.tn.gov', 'www.ccmc.gov', 'payment.ccmc.gov', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'retail.economictimes.indiatimes.com', 'www.hindu.com', 'www.hindu.com', 'www.hinduonnet.com', 'www.resourceinvestor.com', 'www.hindu.com', 'www.thehindu.com', 'indiablooms.com', 'intecexpo.com', 'www.hinduonnet.com', 'articles.timesofindia.indiatimes.com', 'www.hindu.com', 'www.thehindu.com', 'www.thehindubusinessline.com', 'www.hindu.com', 'www.thehindu.com', 'www.thehindubusinessline.com', 'www.hinduonnet.com', 'www.thehindu.com', 'hudku.com', 'timesofindia.indiatimes.com', 'hindu.com', 'www.hindu.com', 'archive.financialexpress.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.hindu.com', 'timesofindia.indiatimes.com', 'www.hindu.com', 'www.livemint.com', 'www.thehindu.com', 'www.iskconhighertaste.com', 'www.bbc.com', 'www.thehindu.com', 'www.deccanherald.com', 'www.hinduonnet.com', 'www.theeyefoundation.com', 'temple.dinamalar.com', 'www.livemint.com', 'timesofindia.indiatimes.com', 'nbnaturepark.com', 'epaper.dailythanthi.com', 'radiomirchi.com', 'www.thehindu.com', 'articles.timesofindia.indiatimes.com', 'books.google.com', 'economictimes.indiatimes.com', 'www.kovaidaily.com', 'economictimes.indiatimes.com', 'siliconindia.com', 'www.thehindu.com', 'www.financialexpress.com', 'articles.economictimes.indiatimes.com', 'sportstaronnet.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehindu.com', 'equitymaster.com', 'www.hindu.com', 'www.hindu.com', 'www.hindu.com', 'www.hindu.com', 'www.hindu.com', 'www.hindu.com', 'www.hinduonnet.com', 'dinakaran.com', 'www.thehindu.com', 'www.thehindubusinessline.com', 'www.thehindu.com', 'eproceedings.worldscinet.com', 'www.thehindu.com', 'www.hindu.com', 'www.hindu.com', 'www.hindu.com', 'articles.economictimes.indiatimes.com', 'www.thehindu.com', 'www.thehindubusinessline.com', 'www.thehindu.com', 'www.hindu.com', 'timesofindia.indiatimes.com', 'www.indiatimes.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.hindu.com', 'www.hinduonnet.com', 'www.hinduonnet.com', 'www.thehindu.com', 'lntecc.com', 'books.google.com', 'www.hindu.com', 'www.thehindu.com', 'news.google.com', 'behindwoods.com', 'www.thehindubusinessline.com', 'indiaprwire.com', 'coimbatoremarathon.com', 'www.hindu.com', 'www.hindu.com', 'timesofindia.indiatimes.com', 'www.hinduonnet.com', 'www.hindu.com', 'www.thehindu.com', 'www.tehelka.com', 'toledoblade.com', 'www.hindu.com', 'books.google.com', 'www.hindu.com', 'epaper.dinamani.com', 'www.thehindu.com', 'www.thehindubusinessline.com', 'www.coimbatore-corporation.com', 'economictimes.indiatimes.com', 'timesofindia.indiatimes.com', 'www.hinduonnet.com', 'books.google.com', 'www.ndtv.com', 'www.hindu.com', 'archive.indianexpress.com', 'www.thehindu.com', 'dinamani.com', 'www.hindu.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.thehindu.com', 'economictimes.indiatimes.com', 'www.newindianexpress.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehindu.com', 'www.hindu.com', 'o3.indiatimes.com', 'hindu.com', 'www.ndtv.com', 'thehindubusinessline.com', 'www.hindu.com', 'www.thehindu.com', 'www.moneycontrol.com', 'www.firstpost.com', 'www.hindu.com', 'www.thehindu.com', 'www.hindu.com', 'www.resourceinvestor.com', 'hudku.com', 'www.hinduonnet.com', 'www.thehindu.com', 'www.hindu.com', 'www.hinduonnet.com', 'www.thehindubusinessline.com', 'www.thehindu.com', 'www.hindu.com', 'www.hinduonnet.com', 'www.hindu.com', 'www.thehindu.com', 'www.thehindu.com', 'www.hindu.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehindu.com', 'www.newindianexpress.com', 'www.thehindu.com', 'www.thehindu.com', 'www.lntidpl.com', 'timesofindia.indiatimes.com', 'www.thehindubusinessline.com', 'www.thehindu.com', 'temple.dinamalar.com', 'dinamalar.com', 'www.thehindu.com', 'www.pppindiadatabase.com', 'www.thehindu.com', 'www.hindu.com', 'www.thehindu.com', 'www.hindu.com', 'indiarailinfo.com', 'www.moneycontrol.com', 'www.hindu.com', 'planetradiocity.com', 'gadgets.ndtv.com', 'www.thehindu.com', 'www.hindu.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehindubusinessline.com', 'citymayors.com', 'www.thehindu.com', 'www.treebo.com', 'timesofindia.indiatimes.com', 'www.hinduonnet.com', 'www.coimbatore-corporation.com', 'economictimes.indiatimes.com', 'www.hindu.com', 'www.thehindu.com', 'www.thehindu.com', 'www.financialexpress.com', 'www.hindu.com', 'articles.timesofindia.indiatimes.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehindubusinessline.com', 'www.hindu.com', 'www.hindu.com', 'www.thehindu.com', 'www.thehindu.com', 'articles.economictimes.indiatimes.com', 'readwhere.com', 'www.hindu.com', 'www.hindu.com', 'www.thehindu.com', 'www.thehindu.com', 'economictimes.indiatimes.com', 'www.thehindu.com', 'www.indiaenvironmentportal.org', 'www.icfre.org', 'afindia.org', 'irfca.org', 'www.sitra.org', 'toledosistercities.org', 'www.nhai.org', ['zoos']]",186096,Require autoconfirmed or confirmed access (no expiry set),176417,21 February 2003,203.199.209.138 ,7749,4,2003-02-21,2003-02,2003
446,446,Tamil Hindu,https://en.wikipedia.org/wiki/Tamil_Hindu,10,2,"['10.1177/006996679903300304', None, None]",[['contributions to indian sociology']],3,0,0,4,0,0,1,0.3,0.0,0.4,0.2,0.0,0.5,1,"['www.thehindu.com', 'www.thehindu.com', 'www.bbc.com', 'food.ndtv.com', 'www.jstor.org', 'tamilnation.org', 'murugan.org', ['contributions to indian sociology']]",53769409,Allow all users (no expiry set),7465,13 April 2017,M.K.Dan ,47,1,2017-04-13,2017-04,2017
447,447,Lahore,https://en.wikipedia.org/wiki/Lahore,210,0,[],[],5,14,0,123,0,1,67,0.023809523809523808,0.06666666666666667,0.5857142857142857,0.0,0.0,0.09047619047619047,0,"['www.pbscensus.gov', 'mail.camara.rj.gov', 'www.pbscensus.gov', 'www.pmd.gov', 'www.pbs.gov', 'www.hko.gov', 'www.nrb.gov', 'www.pbs.gov', 'punjab.gov', 'mail.camara.rj.gov', 'finance.gov', 'lahore.gov', 'www.lahore.gov', 'www.nrb.gov', 'books.google.com', 'books.google.com', 'www.bbc.com', 'www.tribuneindia.com', 'thelahorecity.com', 'books.google.com', 'www.railway-technology.com', 'books.google.com', 'www.milligazette.com', 'homespakistan.com', 'lahore.city-history.com', 'www.gardenvisit.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thenews.com', 'www.ukmediacentre.pwc.com', 'dnd.com', 'www.dawn.com', 'books.google.com', 'books.google.com', 'blogspot.com', 'twitter.com', 'www.storyofpakistan.com', 'pakmet.com', 'dawn.com', 'books.google.com', 'books.google.com', 'tribune.com', 'www.cbsnews.com', 'dawn.com', 'www.dawn.com', 'books.google.com', 'books.google.com', 'lahore.metblogs.com', 'www.expolahore.com', 'www.brecorder.com', 'www.hkttreks.com', 'books.google.com', 'tribune.com', 'www.kroraina.com', 'books.google.com', 'www.lonelyplanet.com', 'lahoreairport.com', 'www.dawn.com', 'books.google.com', 'thenews.com', 'books.google.com', 'books.google.com', 'lahore.city-history.com', 'www.dailytimes.com', 'www.dawn.com', 'books.google.com', 'nation.com', 'www.railjournal.com', 'www.siasat.com', 'christiansinpakistan.com', 'www.dawn.com', 'books.google.com', 'books.google.com', 'arabiclexicon.hawramani.com', 'books.google.com', 'books.google.com', 'www.dawn.com', 'www.thenews.com', 'exoticindiaart.com', 'www.dawn.com', 'nation.com', 'tribune.com', 'books.google.com', 'www.routesonline.com', 'www.economist.com', 'books.google.com', 'www.brecorder.com', 'www.indiatimes.com', 'www.piac.com', 'www.routesonline.com', 'www.dawn.com', 'books.google.com', 'www.dawn.com', 'worldpopulationreview.com', 'www.dailytimes.com', 'www.dailytimes.com', 'books.google.com', 'en.dailypakistan.com', 'tribune.com', 'visitlahore.com', 'books.google.com', 'books.google.com', 'www.thebusinessyear.com', 'thenews.com', 'nation.com', 'www.washingtonpost.com', 'www.routesonline.com', 'www.thenews.com', 'pakvisit.com', 'pakmet.com', 'lahoremarathon.com', 'ghn.globalheritagefund.com', 'www.dailytimes.com', 'tribune.com', 'tribune.com', 'books.google.com', 'books.google.com', 'www.youtube.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.dawn.com', 'tribune.com', 'www.dailytimes.com', 'dailytimes.com', 'www.pakistantoday.com', 'tribune.com', 'www.orientalarchitecture.com', 'www.dawn.com', 'books.google.com', 'dawn.com', 'www.citymayors.com', 'www.ptcl.com', 'www.tribuneindia.com', 'indianexpress.com', 'apnaorg.com', 'whc.unesco.org', 'oic-oci.org', 'www.adb.org', 'www.lahoremetroauraap.org', 'globalsecurity.org']",125315,Allow all users (no expiry set),150710,22 October 2002,204.193.117.66 ,11339,25,2002-10-22,2002-10,2002
448,448,Culture of Iceland,https://en.wikipedia.org/wiki/Culture_of_Iceland,14,1,"['10.1515/fabl.2000.41.1-2.87', None, None]",[['fabula']],0,0,0,4,0,0,9,0.0,0.0,0.2857142857142857,0.07142857142857142,0.0,0.07142857142857142,1,"['www.sciencedaily.com', 'www.einarhakonarson.com', 'www.newyorker.com', 'www.nytimes.com', ['fabula']]",496397,Allow all users (no expiry set),19157,1 March 2004,NuclearWinner ,494,1,2004-03-01,2004-03,2004
449,449,Trabzon,https://en.wikipedia.org/wiki/Trabzon,89,3,"['10.3406/rebyz.1964.1329', '10.4000/eac.1815', '10.5194/hessd-4-439-2007', None, None, None, None, None, None]","[['[[revue des études byzantines'], ['[[études arméniennes contemporaines'], ['hydrology and earth system sciences']]",12,4,0,23,0,0,47,0.1348314606741573,0.0449438202247191,0.25842696629213485,0.033707865168539325,0.0,0.21348314606741572,3,"['trove.nla.gov', 'www.mgm.gov', 'www.mgm.gov', 'www.mgm.gov', 'books.google.com', 'books.google.com', 'ogimet.com', 'books.google.com', 'webcache.googleusercontent.com', 'www.ucuyos.com', 'www.yeniansiklopedi.com', 'www.csmonitor.com', 'www.karalahana.com', 'books.google.com', 'lazuri.com', 'www.weatherbase.com', 'www.ofhayrat.com', 'books.google.com', 'books.google.com', 'karalahana.com', 'www.yeniansiklopedi.com', 'www.nytimes.com', 'books.google.com', 'books.google.com', 'www.thenationalherald.com', 'karalahana.com', 'www.e-bogazici.com', 'www.wdl.org', 'www.wdl.org', 'www.wdl.org', 'www.wdl.org', 'commons.wikimedia.org', 'www.wdl.org', 'www.jstor.org', 'www.jstor.org', 'www.wdl.org', 'islamansiklopedisi.org', 'www.latsis-foundation.org', 'www.wdl.org', ['[[revue des études byzantines'], ['[[études arméniennes contemporaines'], ['hydrology and earth system sciences']]",62653,Allow all users (no expiry set),85780,18 July 2002,216.94.11.2 ,2335,5,2002-07-18,2002-07,2002
450,450,Hazaras,https://en.wikipedia.org/wiki/Hazaras,124,6,"['10.1080/02634939708400997', '10.1126/science.1078311', '10.1371/journal.pone.0034288', '10.1093/molbev/msx177', '10.1371/journal.pone.0161622', '10.1086/383236', None, '12493913', '22470552', '28595347', '27627454', '15077202', None, None, '3314501', None, '5023095', '1181978']","[['central asian survey '], [' science '], ['plos one '], ['molecular biology and evolution'], ['plos one '], ['am. j. hum. genet. ']]",17,4,0,39,0,0,58,0.13709677419354838,0.03225806451612903,0.31451612903225806,0.04838709677419355,0.0,0.21774193548387097,6,"['www.cia.gov', 'www.cia.gov', 'www.loc.gov', 'lcweb2.loc.gov', 'books.google.com', 'books.google.com', 'www.sciencedirect.com', 'www.nbcnews.com', 'www.nytimes.com', 'www.bangkokpost.com', 'pajhwok.com', 'www.nytimes.com', 'www.aljazeera.com', 'nytimes.com', 'tarhenaw.com', 'tribune.com', 'www.csmonitor.com', 'www.tellerreport.com', 'referenceworks.brillonline.com', 'referenceworks.brillonline.com', 'nytimes.com', 'www.nytimes.com', 'hazarapress.com', 'books.google.com', 'ngm.nationalgeographic.com', 'books.google.com', 'www.reuters.com', 'books.google.com', 'www.france24.com', 'dawn.com', 'thediplomat.com', 'www.aljazeera.com', 'books.google.com', 'books.google.com', 'online.wsj.com', 'books.google.com', 'dawn.com', 'www.pdfebooksd.com', 'www.theage.com', 'www.christianitytoday.com', 'referenceworks.brillonline.com', 'www.flickr.com', 'dailytimes.com', 'data.worldbank.org', 'iranicaonline.org', 'www.iranicaonline.org', 'www.cal.org', 'www.bolaq.org', 'iranicaonline.org', 'www.missionfrontiers.org', 'www.jstor.org', 'www.iranicaonline.org', 'iranicaonline.org', 'www.unhcr.org', 'swedishcommittee.org', 'www.jstor.org', 'www.sat7uk.org', 'www.hrw.org', 'www.iranicaonline.org', 'www.washingtoninstitute.org', ['central asian survey '], [' science '], ['plos one '], ['molecular biology and evolution'], ['plos one '], ['am. j. hum. genet. ']]",14131,Require autoconfirmed or confirmed access (no expiry set),76511,25 February 2002,Conversion script ,5288,82,2002-02-25,2002-02,2002
451,451,Como,https://en.wikipedia.org/wiki/Como,33,0,[],[],4,0,0,15,0,0,14,0.12121212121212122,0.0,0.45454545454545453,0.0,0.0,0.12121212121212122,0,"['www.aeroclubcomo.com', 'travel.usnews.com', 'www.comune.com', 'teatrosocialecomo.com', 'meteoblue.com', 'weather-atlas.com', 'www.aeroclubcomo.com', 'www.nytimes.com', 'variety.com', 'answers.com', 'www.ilsole24ore.com', 'www.com', 'www.voyagetips.com', 'books.google.com', 'www.airpullman.com', 'www.npr.org', 'corrosion-doctors.org', 'www.nycgovparks.org', 'openlibrary.org']",60679,Allow all users (no expiry set),37847,6 July 2002,213.45.20.39 ,1061,2,2002-07-06,2002-07,2002
452,452,Louisiana Creole people,https://en.wikipedia.org/wiki/Louisiana_Creole_people,73,0,[],[],7,4,0,20,0,0,42,0.0958904109589041,0.0547945205479452,0.273972602739726,0.0,0.0,0.1506849315068493,0,"['www.nps.gov', 'census.gov', 'www.nps.gov', 'www.nps.gov', 'ebookit.com', 'www.nola.com', 'theneworleanstribune.com', 'avoyelles.com', 'books.google.com', 'iuniverse.com', 'www.katc.com', 'ebookit.com', 'books.google.com', 'www.mylhcv.com', 'www.google.com', 'francolouisiane.com', 'www.everyculture.com', 'www.thenationalherald.com', 'louisianaperspectives.wordpress.com', 'cerebellum1.wordpress.com', 'books.google.com', 'www.lebourdondelalouisiane.com', 'www.louisianacreoledictionary.com', 'www.google.com', 'wcny.org', 'lameca.org', 'www.inmotionaame.org', 'www.knowla.org', 'www.hnoc.org', 'www.zocalopublicsquare.org', 'aaregistry.org']",4167079,Allow all users (no expiry set),78230,23 February 2006,Jorge Stolfi ,2670,10,2006-02-23,2006-02,2006
453,453,Xi'an,https://en.wikipedia.org/wiki/Xi%27an,136,3,"['10.1787/9789264230040-en', '10.1016/j.archoralbio.2011.04.003', None, '21592462', None, None]","[['[[organisation for economic co-operation and development'], ['archives of oral biology']]",4,12,0,66,0,1,50,0.029411764705882353,0.08823529411764706,0.4852941176470588,0.022058823529411766,0.0,0.13970588235294118,2,"['cdc.cma.gov', 'www.xametro.gov', 'www.xa.gov', 'www.edinburgh.gov', 'www.xa.gov', 'www.xatj.gov', 'english.shaanxi.gov', 'www.stats.gov', 'www.edinburgh.gov', 'cdc.cma.gov', 'www.xametro.gov', 'www.xa.gov', 'www.washingtonpost.com', 'www.bbc.com', 'epaper.xiancn.com', 'www.natureindex.com', 'epaper.xiancn.com', 'www.chinadaily.com', 'history.cultural-china.com', 'flyingtiger-cacw.com', 'www.istockanalyst.com', 'chinamuseums.com', 'www.theborneopost.com', 'www.lehmanlaw.com', 'translate.google.com', 'www.chinadaily.com', 'ip138.com', 'english.people.com', 'www.china.com', 'education.yahoo.com', 'books.google.com', 'centreforaviation.com', 'in.reuters.com', 'www.economist.com', 'www.xdz.com', 'gundogar-news.com', 'news.sina.com', 'books.google.com', 'news.xinhuanet.com', 'www.cnbc.com', 'www.huffingtonpost.com', 'www.demographia.com', 'www.britannica.com', 'www.sabahnewstoday.com', 'www.natureindex.com', 'books.google.com', 'www.bestchinanews.com', 'books.google.com', 'books.google.com', 'en.oxforddictionaries.com', 'epaper.xiancn.com', 'english.people.com', 'www.topuniversities.com', 'sg.news.yahoo.com', 'sg.news.yahoo.com', 'www.docin.com', 'books.google.com', 'twins2010.com', 'www.muslim2china.com', 'www.reuters.com', 'www.railwaygazette.com', 'www.huaxia.com', 'newspaperarchive.com', 'www.britannica.com', 'crienglish.com', 'www.usnews.com', 'books.google.com', 'encarta.msn.com', 'www.allroadsleadtochina.com', 'books.google.com', 'china-trade-research.hktdc.com', 'www.collinsdictionary.com', 'www.prnewswire.com', 'science.nationalgeographic.com', 'finance.sina.com', 'www.travelchinaguide.com', 'query.nytimes.com', 'books.google.com', 'china.org', 'www.asiaseia.org', 'www.china.org', 'www.mherrera.org', ['[[organisation for economic co-operation and development'], ['archives of oral biology']]",81263,Allow all users (no expiry set),105395,6 September 2002,Olivier ,3632,23,2002-09-06,2002-09,2002
454,454,Modena,https://en.wikipedia.org/wiki/Modena,15,0,[],[],2,0,0,5,0,0,8,0.13333333333333333,0.0,0.3333333333333333,0.0,0.0,0.13333333333333333,0,"['www.paninigroup.com', 'www.collinsdictionary.com', 'www.com', 'edition.cnn.com', 'beverfood.com', 'visitlakecounty.org', 'en.climate-data.org']",62418,Allow all users (no expiry set),36382,17 July 2002,Gianfranco ,776,1,2002-07-17,2002-07,2002
455,455,Culture of Asia,https://en.wikipedia.org/wiki/Culture_of_Asia,96,5,"['10.1017/s0305741006430241', '10.1016/j.proeng.2016.02.031', '10.1073/pnas.1112743109', '10.1073/pnas.1115430109', '10.3138/utq.29.2.282', None, None, '22645375', '22355109', None, None, None, '3387054', '3309722', None]","[[' the china quarterly ', ' cambridge university press '], ['procedia engineering'], [' proceedings of the national academy of sciences ', ' pnas '], [' proceedings of the national academy of sciences', 'pnas'], ['university of toronto quarterly']]",23,3,0,35,0,0,30,0.23958333333333334,0.03125,0.3645833333333333,0.052083333333333336,0.0,0.3229166666666667,5,"['www.nla.gov', 'e-reports-ext.llnl.gov', 'www.loc.gov', 'www.thoughtco.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'books.google.com', 'dimensionsofculture.com', 'www.britannica.com', 'books.google.com', 'www.britannica.com', 'www.ricearoni.com', 'books.google.com', 'books.google.com', 'thediplomat.com', 'books.google.com', 'www.dimensionsofculture.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'www.britannica.com', 'www.amitavacharya.com', 'books.google.com', 'books.google.com', 'www.allempires.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.omniglot.com', 'history.intellichristian.com', 'books.google.com', 'www.britannica.com', 'www.realcleardefense.com', 'asiasociety.org', 'www.jewishvirtuallibrary.org', 'www.pewforum.org', 'www.worldcat.org', 'www.pewforum.org', 'web-japan.org', 'asiasociety.org', 'asiasociety.org', 'unstats.un.org', 'www.pewforum.org', 'asiasociety.org', 'www.pewforum.org', 'whc.unesco.org', 'www.nationalgeographic.org', 'www.fpmtmongolia.org', 'www.pewforum.org', 'assets.pewresearch.org', 'npr.org', 'www.un.org', 'www.pewforum.org', 'www.pewforum.org', 'www.pewforum.org', 'www.pewforum.org', [' the china quarterly ', ' cambridge university press '], ['procedia engineering'], [' proceedings of the national academy of sciences ', ' pnas '], [' proceedings of the national academy of sciences', 'pnas'], ['university of toronto quarterly']]",1738605,Allow all users (no expiry set),99107,14 April 2005,220.226.30.178 ,2103,6,2005-04-14,2005-04,2005
456,456,Culture of England,https://en.wikipedia.org/wiki/Culture_of_England,450,8,"['10.2307/898796', '10.1038/1811754a0', '10.18111/9789284421152', '10.1017/cbo9781139097192', '10.5040/9781472575692', '10.1017/cbo9780511819520', '10.2307/2595542', None, None, None, None, None, None, None, None, None, None, None, None, None, None]","[['notes'], ['nature'], ['world tourism organization '], [' [[cambridge university press'], [' [[bloomsbury publishing'], [' [[cambridge university press'], ['the economic history review']]",38,16,0,90,0,17,281,0.08444444444444445,0.035555555555555556,0.2,0.017777777777777778,0.0,0.13777777777777778,7,"['www.gov', 'number10.gov', 'www.gov', 'www.gov', 'www.gov', 'www.gov', 'www.gov', 'www.cambridge.gov', 'www.gov', 'www.nationalarchives.gov', 'www.gov', 'www.gov', 'www.cambridge.gov', 'www.insolvency.gov', 'www.gov', 'www.legislation.gov', 'www.ealingstudios.com', 'www.sportinglife.com', 'www.historic-uk.com', 'projectbritain.com', 'www.artinfo.com', 'www.travour.com', 'books.google.com', 'www.cricinfo.com', 'yourdictionary.com', 'www.nytimes.com', 'www.redorbit.com', 'www.timescolonist.com', 'www.englishbreakfastsociety.com', 'www.britannica.com', 'www.thoughtco.com', 'www.whatdadcooked.com', 'fifa.com', 'www.all-about-afternoon-tea.com', 'www.tripsavvy.com', 'www.pgatour.com', 'thedrinksbusiness.com', 'ratetea.com', 'www.economist.com', 'www.bbc.com', 'www.waitrose.com', 'statisticalyearbook11.ry.com', 'www.cheese.com', 'www.time.com', 'beerandbrewing.com', 'ebert.com', 'www.topuniversities.com', 'books.google.com', 'www.cheese.com', 'www.britannica.com', 'uk.encarta.msn.com', 'books.google.com', 'www.cricinfo.com', 'books.google.com', 'www.gordonramsayrestaurants.com', 'chilliandmint.com', 'www.channel4.com', 'www.britannica.com', 'www.timeshighereducation.com', 'www.economist.com', 'www.anyoneforpimms.com', 'www.britannica.com', 'www.theworlds50best.com', 'www.tennisfame.com', 'projectbritain.com', 'drinks.seriouseats.com', 'www.itv.com', 'www.bbc.com', 'www.lonelyplanet.com', 'www.all-about-afternoon-tea.com', 'www.dezeen.com', 'everynoise.com', 'longleyfarm.com', 'www.historytoday.com', 'edition.cnn.com', 'coventmarket.com', 'www.beeradvocate.com', 'rankings.ft.com', 'drinkstack.com', 'www.beeradvocate.com', 'rugbyfootballhistory.com', 'www.timeshighereducation.com', 'history.com', 'www.cheese.com', 'www.nytimes.com', 'www.britannica.com', 'dictionary.law.com', 'books.google.com', 'www.bbc.com', 'www.ppluk.com', 'www.britannica.com', 'britishfoodhistory.com', 'bleacherreport.com', 'uk.encarta.msn.com', 'lovefood.com', 'greatbritishmeat.com', 'www.englandanthem.com', 'encarta.msn.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'www.bartleby.com', 'slate.com', 'www.americanheritage.com', 'www.uhy-uk.com', 'www.essentially-england.com', 'www.english-heritage.org', 'www.english-heritage.org', 'www.artscouncil.org', 'www.neoda.org', 'www.tate.org', 'visitbritain.org', 'rts.org', 'rsliterature.org', 'cccbr.org', 'www.rhs.org', 'www.english-heritage.org', 'www.thersa.org', 'www.bfi.org', 'royalsociety.org', 'www.sustainweb.org', 'www.camra.org', 'www.britishmuseum.org', 'www.foodtimeline.org', 'www.roh.org', 'smarthistory.org', 'www.camra.org', 'abbey.org', 'www.stone-circles.org', 'www.socialisteducation.org', 'blog.english-heritage.org', 'www.campaignforrealfarming.org', 'royalsociety.org', 'royalsociety.org', 'www.tate.org', 'www.sweca.org', 'www.ihbc.org', 'www.seafish.org', 'www.ofcom.org', 'www.metmuseum.org', 'www.english-heritage.org', 'shop.ashmolean.org', 'piers.org', 'historicengland.org', ['notes'], ['nature'], ['world tourism organization '], [' [[cambridge university press'], [' [[bloomsbury publishing'], [' [[cambridge university press'], ['the economic history review']]",60603911,Allow all users (no expiry set),239191,18 November 2004,Thewayforward ,3839,3,2004-11-18,2004-11,2004
457,457,Dortmund,https://en.wikipedia.org/wiki/Dortmund,99,0,[],[],5,0,0,13,0,0,81,0.050505050505050504,0.0,0.13131313131313133,0.0,0.0,0.050505050505050504,0,"['www.natureindex.com', 'www.aerotelegraph.com', 'www.innovation-cities.com', 'frankfurt-expat.com', 'www.cbsnews.com', 'www.musicbusinessworldwide.com', 'thebeergeek.com', 'www.mhp.com', 'digitalhublogistics.com', 'www.nytimes.com', 'botschaft-konsulat.com', 'www.tripadvisor.com', 'edition.cnn.com', 'www.bitkom.org', 'www.ibo.org', 'backtonormandy.org', 'www.lwl.org', 'www.kirchentag.org']",149349,Allow all users (no expiry set),121715,20 November 2002,WojPob ,1687,4,2002-11-20,2002-11,2002
458,458,Pomerania,https://en.wikipedia.org/wiki/Pomerania,46,0,[],[],1,0,0,5,0,0,40,0.021739130434782608,0.0,0.10869565217391304,0.0,0.0,0.021739130434782608,0,"['www.bartleby.com', 'books.google.com', 'books.google.com', 'www.bartleby.com', 'www.britannica.com', 'midiacidada.org']",24261,Allow all users (no expiry set),47015,2 October 2001,MichaelTinkler ,1563,1,2001-10-02,2001-10,2001
459,459,Ancient Macedonians,https://en.wikipedia.org/wiki/Ancient_Macedonians,445,6,"['10.1515/9783110532135', '10.1515/9783110532135-013', '10.12681/bgsg.17141', '10.1111/1468-0092.00106', '10.1093/cq/53.2.510', '10.3765/bls.v25i1.1180', None, None, None, None, None, None, None, None, None, None, None, None]","[['de gruyter'], ['[[de gruyter'], ['bulletin of the geological society of greece', 'proceedings of the 11th international congress'], ['oxford journal of archaeology'], ['the classical quarterly'], [' annual meeting of the berkeley linguistics society']]",4,0,0,101,0,0,334,0.008988764044943821,0.0,0.22696629213483147,0.01348314606741573,0.0,0.02247191011235955,6,"['books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.seeker.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'gradworks.umi.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'greece.greekreporter.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.oxforddictionaries.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.gutenberg.org', 'macedonia-evidence.org', 'www.livius.org', 'macedonia-evidence.org', ['de gruyter'], ['[[de gruyter'], ['bulletin of the geological society of greece', 'proceedings of the 11th international congress'], ['oxford journal of archaeology'], ['the classical quarterly'], [' annual meeting of the berkeley linguistics society']]",2417624,Require administrator access (no expiry set),176392,10 August 2005,Alex '05 ,3043,0,2005-08-10,2005-08,2005
460,460,Sicilians,https://en.wikipedia.org/wiki/Sicilians,123,29,"['10.3764/aja.115.3.0447', '10.1038/ejhg.2015.124', '10.1371/journal.pone.0192269', '10.6092/2037-4488/1940', '10.1038/ejhg.2008.120', '10.1163/1570058982641743', '10.1038/ejhg.2015.233', '10.1038/ejhg.2017.18', '10.3390/geosciences8070253', '10.1016/j.ajhg.2008.10.012', '10.1186/s12863-015-0293-x', '10.1371/journal.pone.0096074', '10.1111/j.1529-8817.2005.00224.x', '10.1371/journal.pone.0050794', '10.6092/2037-4488/1942', '10.1038/s41598-017-01802-4', '10.1073/pnas.1320811111', '10.1590/s1415-47572004000200002', '10.1002/ajpa.10265', '10.1111/j.1469-1809.2007.00414.x', '10.1038/ejhg.2008.258', '10.1371/journal.pone.0043759', '10.1126/sciadv.aaw3492', '10.1111/ahg.12328', '10.1038/srep32513', '10.1098/rspb.2019.0471', '10.1038/s41431-019-0466-6', None, '26173964', '29522542', None, '18685561', None, '26554880', '28272534', None, '18976729', '26553317', '24788788', '16626331', '23251386', None, '28512355', '24927591', None, '12772214', '18269686', '19156170', '22984441', '31517044', '31192450', '27582244', '31039721', '31285530', None, '4757772', '5844529', None, '2985948', None, '5070887', '5437898', None, '2668035', '4640365', '4005757', None, '3519480', None, '5434004', '4078858', None, None, None, '2947089', '3440425', '6726452', '6851683', '5007512', '6532504', '6871633']","[['american journal of archaeology'], ['european journal of human genetics '], ['plos one'], ['aristonothos 4 '], ['european journal of human genetics'], ['arabica'], ['european journal of human genetics '], ['european journal of human genetics '], ['geosciences '], ['the american journal of human genetics'], ['bmc genetics'], ['plos one '], ['annals of human genetics '], ['plos one'], ['aristonothos 4 '], ['scientific reports '], ['proceedings of the national academy of sciences of the united states of america '], ['genetics and molecular biology '], [' american journal of physical anthropology'], ['annals of human genetics '], [' european journal of human genetics'], ['plos one '], ['science advances '], ['annals of human genetics '], [' nature'], ['proceedings of the royal society b'], ['european journal of human genetics ']]",6,0,0,27,0,0,61,0.04878048780487805,0.0,0.21951219512195122,0.23577235772357724,0.0,0.2845528455284553,27,"['www.ancientlibrary.com', 'books.google.com', 'siciliangodmother.com', 'books.google.com', 'books.google.com', 'www.thethinkingtraveller.com', 'www.bestofsicily.com', 'www.experiencefestival.com', 'referenceworks.brillonline.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.italymagazine.com', 'books.google.com', 'experiencesicily.com', 'books.google.com', 'www.haaretz.com', 'www.businesstimes.com', 'books.google.com', 'theculturetrip.com', 'www.haaretz.com', 'books.google.com', 'www.timesofsicily.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.gatestoneinstitute.org', 'linguistlist.org', 'www.michaelfreund.org', 'www.newadvent.org', 'whc.unesco.org', 'www.usefinternational.org', ['american journal of archaeology'], ['european journal of human genetics '], ['plos one'], ['aristonothos 4 '], ['european journal of human genetics'], ['arabica'], ['european journal of human genetics '], ['european journal of human genetics '], ['geosciences '], ['the american journal of human genetics'], ['bmc genetics'], ['plos one '], ['annals of human genetics '], ['plos one'], ['aristonothos 4 '], ['scientific reports '], ['proceedings of the national academy of sciences of the united states of america '], ['genetics and molecular biology '], [' american journal of physical anthropology'], ['annals of human genetics '], [' european journal of human genetics'], ['plos one '], ['science advances '], ['annals of human genetics '], [' nature'], ['proceedings of the royal society b'], ['european journal of human genetics ']]",1070829,Allow all users (no expiry set),94789,15 October 2004,68.157.156.180 ,1207,8,2004-10-15,2004-10,2004
461,461,Creuse,https://en.wikipedia.org/wiki/Creuse,5,0,[],[],0,0,0,2,0,0,3,0.0,0.0,0.4,0.0,0.0,0.0,0,"['www.encreuse.com', 'www.jedecouvrelafrance.com']",90551,Allow all users (no expiry set),20938,24 September 2002,Olivier ,355,10,2002-09-24,2002-09,2002
462,462,Lingnan culture,https://en.wikipedia.org/wiki/Lingnan_culture,53,2,"['10.1016/j.jep.2019.112491', None, None]",[['journal of ethnopharmacology ']],2,2,0,18,0,0,29,0.03773584905660377,0.03773584905660377,0.33962264150943394,0.03773584905660377,0.0,0.11320754716981132,1,"['catalogue.nla.gov', 'www.lcsd.gov', 'read01.com', 'lulu.com', 'read01.com', 'www.chinanews.com', 'thefadingfolkmemory.weebly.com', 'www.atoomu.com', 'hk.crntt.com', 'read01.com', 'www.gdwh.com', 'www.scmp.com', 'www.chinabaike.com', 'lulu.com', 'read01.com', 'www.cantoneseculture.com', 'read01.com', 'news.sina.com', 'www.chinatyxk.com', 'read01.com', 'en.unesco.org', 'www.huayuqiao.org', ['journal of ethnopharmacology ']]",2042987,Allow all users (no expiry set),68320,14 June 2005,Dpr ,860,3,2005-06-14,2005-06,2005
463,463,Bilbao,https://en.wikipedia.org/wiki/Bilbao,193,0,[],[],7,0,0,62,0,0,124,0.03626943005181347,0.0,0.32124352331606215,0.0,0.0,0.03626943005181347,0,"['www.elcorreo.com', 'www.worldmayor.com', 'www.periodistasvascos.com', 'www.asierpolo.com', 'www.deia.com', 'soccernet.espn.go.com', 'moovitapp.com', 'population-statistics.com', 'www.elcorreo.com', 'www.elcorreo.com', 'euskonews.com', 'www.periodistasvascos.com', 'www.periodistasvascos.com', 'www.lavanguardia.com', 'www.alhondigabilbao.com', 'www.periodistasvascos.com', 'www.deia.com', 'www.elcorreo.com', 'www.elcorreo.com', 'bajoelagua.com', 'bilbaohiria.com', 'www.deia.com', 'www.worldmayor.com', 'moovitapp.com', 'www.elcorreo.com', 'www.elcorreodigital.com', 'www.collinsdictionary.com', 'www.periodistasvascos.com', 'www.elcorreo.com', 'www.elcorreo.com', 'www.vanityfair.com', 'www.elcorreo.com', 'www.periodistasvascos.com', 'athletic-zurekin.com', 'www.deia.com', 'www.alhondigabilbao.com', 'www.elcorreodigital.com', 'www.periodistasvascos.com', 'www.museobilbao.com', 'www.elcorreo.com', 'elviajero.elpais.com', 'www.periodistasvascos.com', 'www.elcorreodigital.com', 'www.elcorreo.com', 'www2.deia.com', 'books.google.com', 'www.elpais.com', 'bilbaobasket.elcorreo.com', 'ogimet.com', 'servicios.elcorreodigital.com', 'euskonews.com', 'descargas.cervantesvirtual.com', 'info.elcorreo.com', 'www.elcorreo.com', 'www.proyectosbilbao.com', 'www.periodistasvascos.com', 'www.deia.com', 'www.elpais.com', 'www.leekuanyewworldcityprize.com', 'footballcitizens.com', 'en.oxforddictionaries.com', 'euskonews.com', 'en.unesco.org', 'www.bilbaoria2000.org', 'en.unesco.org', 'unesdoc.unesco.org', 'www.euskal-museoa.org', 'euskomedia.org', 'euskomedia.org']",68029,Allow all users (no expiry set),161010,5 August 2002,207.253.140.103 ,2409,7,2002-08-05,2002-08,2002
464,464,Minangkabau culture,https://en.wikipedia.org/wiki/Minangkabau_culture,18,2,"['10.1046/j.1440-6047.2001.00201.x', '10.1353/atj.2003.0025', '11708602', None, None, None]","[['asia pacific journal of clinical nutrition ', 'blackwell synergy '], ['asian theatre journal ']]",0,1,0,7,0,0,8,0.0,0.05555555555555555,0.3888888888888889,0.1111111111111111,0.0,0.16666666666666666,2,"['lcweb2.loc.gov', 'www.bbc.com', 'www.cnngo.com', 'www.thejakartapost.com', 'theconversation.com', 'www.cnngo.com', 'kompas.com', 'www.thejakartapost.com', ['asia pacific journal of clinical nutrition ', 'blackwell synergy '], ['asian theatre journal ']]",66075231,Allow all users (no expiry set),26680,11 December 2020,Xcelltrasi ,58,0,2020-12-11,2020-12,2020
465,465,Arrifana (Aljezur),https://en.wikipedia.org/wiki/Arrifana_(Aljezur),28,0,[],[],0,0,0,11,0,0,17,0.0,0.0,0.39285714285714285,0.0,0.0,0.0,0,"['www.iberian-escapes.com', 'rotavicentina.com', 'thesurfatlas.com', 'www.businessinsider.com', 'algarvedailynews.com', 'www.iberian-escapes.com', 'www.vice.com', 'culturanoporto.canalblog.com', 'surfergalaxy.com', 'blog.algarveholidaylets.com', 'rotavicentina.com']",5313902,Allow all users (no expiry set),16194,27 May 2006,Timkevan ,25,0,2006-05-27,2006-05,2006
466,466,Culture of Azerbaijan,https://en.wikipedia.org/wiki/Culture_of_Azerbaijan,65,0,[],[],6,2,0,23,0,0,34,0.09230769230769231,0.03076923076923077,0.35384615384615387,0.0,0.0,0.12307692307692308,0,"['lcweb2.loc.gov', 'mfa.gov', 'www.washingtonpost.com', 'www.britannica.com', 'www.britannica.com', 'www.azer.com', 'www.azer.com', 'www.echo-az.com', 'azerembsof.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'bangkokcompanies.com', 'everyculture.com', 'www.wtmlondon.com', 'www.iranica.com', 'books.google.com', 'www.hauntedink.com', 'hankooki.com', 'azeriyoungsters.blogspot.com', 'www.nytimes.com', 'books.google.com', 'anspress.com', 'everyculture.com', 'books.google.com', 'ich.unesco.org', 'features.pewforum.org', 'isesco.org', 'eurasianet.org', 'azerembassy-kuwait.org', 'www.isesco.org']",2071240,Allow all users (no expiry set),53175,19 June 2005,Dpr ,569,0,2005-06-19,2005-06,2005
467,467,Corsica,https://en.wikipedia.org/wiki/Corsica,72,0,[],[],4,1,0,17,0,2,48,0.05555555555555555,0.013888888888888888,0.2361111111111111,0.0,0.0,0.06944444444444445,0,"['www.weather.gov', 'www.corsica-isula.com', 'www.economist.com', 'articles.baltimoresun.com', 'www.mobylines.com', 'tempsreel.nouvelobs.com', 'www.corsicaexperience.com', 'www.rue89.com', 'books.google.com', 'french-at-a-touch.com', 'globaltwitcher.com', 'books.google.com', 'www.cnn.com', 'arthursclassicnovels.com', 'www.nytimes.com', 'www.corsica-isula.com', 'yellowbordermagazine.com', 'www.meteofrance.com', 'glottolog.org', 'www.unesco.org', 'wayback.archive-it.org', 'www.prehistoire-corse.org']",5714828,Allow all users (no expiry set),76539,4 December 2001,209.232.151.xxx ,2888,11,2001-12-04,2001-12,2001
468,468,Prekmurje,https://en.wikipedia.org/wiki/Prekmurje,8,0,[],[],0,0,0,0,0,0,8,0.0,0.0,0.0,0.0,0.0,0.0,0,[],983371,Allow all users (no expiry set),19183,14 September 2004,193.77.157.91 ,454,1,2004-09-14,2004-09,2004
469,469,Aosta Valley,https://en.wikipedia.org/wiki/Aosta_Valley,42,2,"['10.2307/40142443', '10.1080/01434632.1984.9994177', None, None, None, None]","[['world literature today '], ['journal of multilingual and multicultural development ']]",6,0,0,3,0,0,31,0.14285714285714285,0.0,0.07142857142857142,0.047619047619047616,0.0,0.19047619047619047,2,"['books.google.com', 'valdostadailytimes.com', 'books.google.com', 'www.heraldica.org', 'www.fondchanoux.org', 'www.fondchanoux.org', 'hdi.globaldatalab.org', 'eso.org', 'www.fondchanoux.org', ['world literature today '], ['journal of multilingual and multicultural development ']]",301306,Allow all users (no expiry set),30563,21 August 2003,Pietro ,993,1,2003-08-21,2003-08,2003
470,470,Dera Ismail Khan District,https://en.wikipedia.org/wiki/Dera_Ismail_Khan_District,14,0,[],[],2,6,0,3,0,0,3,0.14285714285714285,0.42857142857142855,0.21428571428571427,0.0,0.0,0.5714285714285714,0,"['dikhan.kp.gov', 'www.nrb.gov', 'pk.usembassy.gov', 'www.pbs.gov', 'www.pbscensus.gov', 'www.panwfp.gov', 'books.google.com', 'www.google.com', 'www.britannica.com', 'waseb.org', 'www.jstor.org']",988585,Allow all users (no expiry set),18844,15 September 2004,65.195.62.33 ,758,3,2004-09-15,2004-09,2004
471,471,Tang dynasty,https://en.wikipedia.org/wiki/Tang_dynasty,44,1,"['10.1111/0020-8833.00053', None, None]",[[' [[international studies quarterly']],3,0,0,15,0,0,25,0.06818181818181818,0.0,0.3409090909090909,0.022727272727272728,0.0,0.09090909090909091,1,"['books.google.com', 'books.google.com', 'www.dictionary.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'referenceworks.brillonline.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'artsbma.org', 'artsbma.org', 'thetangdynasty.org', [' [[international studies quarterly']]",43455,Allow all users (no expiry set),168658,9 March 2002,63.192.137.21 ,7385,11,2002-03-09,2002-03,2002
472,472,Frogs in culture,https://en.wikipedia.org/wiki/Frogs_in_culture,42,0,[],[],6,0,0,12,0,1,23,0.14285714285714285,0.0,0.2857142857142857,0.0,0.0,0.14285714285714285,0,"['articles.timesofindia.indiatimes.com', 'www.imdb.com', 'www.smh.com', 'www.bogleech.com', 'tv.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.fastcompany.com', 'www.bogleech.com', 'time.com', 'ctext.org', 'www.jstor.org', 'www.the-leaky-cauldron.org', 'tropes.org', 'www.nationalgallery.org', 'www.bopsecrets.org']",3865065,Allow all users (no expiry set),24305,27 January 2006,Samsara ,627,1,2006-01-27,2006-01,2006
473,473,Mersin,https://en.wikipedia.org/wiki/Mersin,20,0,[],[],3,4,0,6,0,0,7,0.15,0.2,0.3,0.0,0.0,0.35,0,"['www.mersin2013.gov', 'www.mersin2013.gov', 'www.mersin.gov', 'www.mgm.gov', 'www.zaman.com', 'www.hurriyetdailynews.com', 'www.forummersin.com', 'www.haberturk.com', 'www.nufusu.com', 'en.firatnews.com', 'www.wdl.org', 'www.wdl.org', 'www.wdl.org']",1146241,Allow all users (no expiry set),32277,8 November 2004,Leandros ,1117,4,2004-11-08,2004-11,2004
474,474,Culture of Albania,https://en.wikipedia.org/wiki/Culture_of_Albania,67,0,[],[],12,0,0,28,0,0,27,0.1791044776119403,0.0,0.417910447761194,0.0,0.0,0.1791044776119403,0,"['books.google.com', 'books.google.com', 'bbc.com', 'books.google.com', 'books.google.com', 'apnews.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'shqiptarja.com', 'books.google.com', 'books.google.com', 'books.google.com', 'ijoer.com', 'ynetnews.com', 'books.google.com', 'www.lesartsturcs.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.balkaninsight.com', 'books.google.com', 'books.google.com', 'books.google.com', 'gazetaexpress.com', 'books.google.com', 'www.jewishvirtuallibrary.org', 'ich.unesco.org', 'frosina.org', 'whc.unesco.org', 'unesco.org', 'unesco.org', 'whc.unesco.org', 'mirror.undp.org', 'yadvashem.org', 'eastagri.org', 'biblicalstudies.org', 'www.jewishvirtuallibrary.org']",167218,Allow all users (no expiry set),62290,9 January 2003,Dori ,609,5,2003-01-09,2003-01,2003
475,475,Lika,https://en.wikipedia.org/wiki/Lika,15,0,[],[],2,0,0,3,0,0,10,0.13333333333333333,0.0,0.2,0.0,0.0,0.13333333333333333,0,"['lika-gastro.com', 'books.google.com', 'lika-gastro.com', 'www.cambridge.org', 'ia360925.us.archive.org']",449899,Allow all users (no expiry set),20153,1 February 2004,Igor~enwiki ,723,0,2004-02-01,2004-02,2004
476,476,Larnaca,https://en.wikipedia.org/wiki/Larnaca,14,0,[],[],2,4,0,0,0,0,8,0.14285714285714285,0.2857142857142857,0.0,0.0,0.0,0.42857142857142855,0,"['www.mof.gov', 'www.mfa.gov', 'www.moa.gov', 'www.cystat.gov', 'www.larnaka.org', 'meteo-climat-bzh.dyndns.org']",287852,Allow all users (no expiry set),26234,4 August 2003,194.219.160.131 ,1299,2,2003-08-04,2003-08,2003
477,477,Saurashtra people,https://en.wikipedia.org/wiki/Saurashtra_people,84,1,"['10.1017/s0035869x00099020', None, None]",[['journal of the royal asiatic society']],2,0,0,67,0,1,13,0.023809523809523808,0.0,0.7976190476190477,0.011904761904761904,0.0,0.03571428571428571,1,"['www.hindustantimes.com', 'www.thehindu.com', 'books.google.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.boloji.com', 'books.google.com', 'www.thebetterindia.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.thehindu.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'rjisacjournal.com', 'www.newindianexpress.com', 'www.thehindu.com', 'www.popsci.com', 'www.deccanchronicle.com', 'www.thehindu.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'books.google.com', 'food.ndtv.com', 'books.google.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'www.telegraphindia.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'www.ethnologue.com', 'www.boloji.com', 'www.thehindu.com', 'food.manoramaonline.com', 'www.indulgexpress.com', 'www.indiapost.com', 'www.thehindu.com', 'books.google.com', 'www.deccanchronicle.com', 'books.google.com', 'www.vepachedu.org', 'indiadivine.org', ['journal of the royal asiatic society']]",29247800,Allow all users (no expiry set),56438,18 October 2010,Shabdarth ,1065,44,2010-10-18,2010-10,2010
478,478,Aromanians,https://en.wikipedia.org/wiki/Aromanians,79,4,"['10.1038/ejhg.2010.146', '10.1215/10474552-15-4-115', '10.1111/j.1469-1809.2005.00251.x', '10.17951/rh.2016.41.213', '20736979', None, '16759179', None, '3039512', None, None, None]","[['european journal of human genetics'], ['mediterranean quarterly'], [' annals of human genetics '], ['res historica ']]",9,4,0,21,0,0,41,0.11392405063291139,0.05063291139240506,0.26582278481012656,0.05063291139240506,0.0,0.21518987341772153,4,"['www.stat.gov', 'www.popis.gov', 'webrzs.stat.gov', 'www.instat.gov', 'britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'search.proquest.com', 'search.proquest.com', 'books.google.com', 'bjuniornewblog.blogspot.com', 'books.google.com', 'www.ceeol.com', 'es.scribd.com', 'books.google.com', 'www.ceeol.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'vatopaidi.wordpress.com', 'books.google.com', 'eblul.org', 'eblul.org', 'cincari.org', 'escholarship.org', 'www.semanticscholar.org', 'www.eurominority.org', 'books.openedition.org', 'www.farsarotul.org', 'etar.org', ['european journal of human genetics'], ['mediterranean quarterly'], [' annals of human genetics '], ['res historica ']]",323104,Allow all users (no expiry set),76181,20 September 2003,Bogdangiusca ,4684,6,2003-09-20,2003-09,2003
479,479,Dakshina Kannada,https://en.wikipedia.org/wiki/Dakshina_Kannada,139,2,"['10.6024/jmbai.2013.55.2.01768-07', '10.1136/tobaccocontrol-2013-051404', None, '24789606', None, None]","[['marine biological association of india', 'journal of the marine biological association of india'], ['tobacco control']]",10,10,0,80,0,0,37,0.07194244604316546,0.07194244604316546,0.5755395683453237,0.014388489208633094,0.0,0.15827338129496402,2,"['www.censusindia.gov', 'dspace.wbpublibnet.gov', 'imdpune.gov', 'www.cpcri.gov', 'www.kpwd.gov', 'gcmd.nasa.gov', 'censusindia.gov', 'www.cia.gov', 'cgwb.gov', 'imdpune.gov', 'news.nationalpost.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.daijiworld.com', 'timesofindia.indiatimes.com', 'www.thehindubusinessline.com', 'rediff.com', 'weather-and-climate.com', 'books.google.com', 'pppinindia.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehindu.com', 'www.deccanherald.com', 'books.google.com', 'www.thehindu.com', 'articles.timesofindia.indiatimes.com', 'www.thehindubusinessline.com', 'www.arvindguptatoys.com', 'www.hindu.com', 'timesofindia.indiatimes.com', 'www.thehindubusinessline.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'www.newindianexpress.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehindu.com', 'economictimes.indiatimes.com', 'www.thehindu.com', 'www.icicihfc.com', 'www.thehindu.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.daijiworld.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehindu.com', 'www.newindianexpress.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.thehindu.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'www.hindu.com', 'www.thehindu.com', 'www.deccanherald.com', 'www.hindu.com', 'www.deccanchronicle.com', 'www.firstpost.com', 'books.google.com', 'books.google.com', 'www.karnataka.com', 'www.thehindu.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.daijiworld.com', 'mangalorean.com', 'books.google.com', 'www.hindu.com', 'www.hindu.com', 'www.daijiworld.com', 'elevation.maplogs.com', 'indianhistorybooks.files.wordpress.com', 'www.deccanherald.com', 'www.newmangalore-port.com', 'www.livemint.com', 'www.daftlogic.com', 'www.daijiworld.com', 'www.deccanherald.com', 'www.daijiworld.com', 'www.fallingrain.com', 'www.khaleejtimes.com', 'karnataka.com', 'timesofindia.indiatimes.com', 'provglo.org', 'www.unep.org', 'www.nhai.org', 'www.cofmangalore.org', 'climate-data.org', 'www.jstor.org', 'www.commonlii.org', 'www.campco.org', 'climate-data.org', 'www.sobiad.org', ['marine biological association of india', 'journal of the marine biological association of india'], ['tobacco control']]",883452,Allow all users (no expiry set),87576,7 August 2004,Tom Radulovich ,2026,6,2004-08-07,2004-08,2004
480,480,Madheshi people,https://en.wikipedia.org/wiki/Madheshi_people,54,6,"['10.1080/09700161.2011.576099', '10.1111/j.1749-8171.2011.00314.x', '10.1111/1467-9655.13025', '10.1080/03068374.2014.909627', '10.1017/s0026749x15000438', '10.1080/02666958108715821', None, None, None, None, None, None, None, None, None, None, None, None]","[['strategic analysis '], ['religion compass '], ['journal of the royal anthropological institute '], ['asian affairs '], ['modern asian studies '], ['journal of muslim minority affairs ']]",8,1,0,15,0,0,24,0.14814814814814814,0.018518518518518517,0.2777777777777778,0.1111111111111111,0.0,0.2777777777777778,6,"['www.loc.gov', 'nepalitimes.com', 'madhesh.com', 'www.ashraya-nepal.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'thediplomat.com', 'www.bbc.com', 'nepalitimes.com', 'books.google.com', 'www.aljazeera.com', 'books.google.com', 'books.google.com', 'indianexpress.com', 'coin.fao.org', 'unstats.un.org', 'lib.icimod.org', 'www.satp.org', 'unpo.org', 'apjcn.nhri.org', 'cscenter.org', 'fwld.org', ['strategic analysis '], ['religion compass '], ['journal of the royal anthropological institute '], ['asian affairs '], ['modern asian studies '], ['journal of muslim minority affairs ']]",8062531,Require autoconfirmed or confirmed access (no expiry set),30386,22 November 2006,Dryman ,1829,0,2006-11-22,2006-11,2006
481,481,Nakhchivan (city),https://en.wikipedia.org/wiki/Nakhchivan_(city),81,0,[],[],6,5,0,12,0,0,58,0.07407407407407407,0.06172839506172839,0.14814814814814814,0.0,0.0,0.13580246913580246,0,"['ftp.atdd.noaa.gov', 'www.stat.gov', 'www.mincom.gov', 'stat.gov', 'www.meclis.gov', 'uefa.com', 'uefa.com', 'www.dw.com', 'azerifootball.com', 'www.bbc.com', 'library.untraveledroad.com', 'www.noahsarksearch.com', 'nakhchivan2014.com', 'www.fni.com', 'capital.trendaz.com', 'www.ekhokavkaza.com', 'transit.parovoz.com', 'www.belediyye.org', 'whc.unesco.org', 'unesco.org', 'www.iranicaonline.org', 'www.iranicaonline.org', 'www.iranicaonline.org']",1492960,Allow all users (no expiry set),46916,11 February 2005,Golbez ,864,0,2005-02-11,2005-02,2005
482,482,Kumaoni people,https://en.wikipedia.org/wiki/Kumaoni_people,18,1,"['10.2307/600927', None, None]",[['journal of the american oriental society']],3,1,0,9,0,0,4,0.16666666666666666,0.05555555555555555,0.5,0.05555555555555555,0.0,0.2777777777777778,1,"['censusindia.gov', 'euttaranchal.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'tribuneindia.com', 'www.jagran.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.iloveindia.com', 'www.unesco.org', 'www.himalayanlanguages.org', 'www.unesco.org', ['journal of the american oriental society']]",22531422,Allow all users (no expiry set),13578,23 April 2009,Kalikumaun ,1441,2,2009-04-23,2009-04,2009
483,483,Mappila Muslims,https://en.wikipedia.org/wiki/Mappila_Muslims,80,3,"['10.33306/mjssh/31', None, None]",[['muallim journal of social sciences and humanities']],2,4,0,40,0,0,31,0.025,0.05,0.5,0.0375,0.0,0.1125,1,"['www.keralapsc.gov', 'censusindia.gov', 'www.censusindia.gov', 'kerala.gov', 'books.google.com', 'books.google.com', 'traveller.outlookindia.com', 'www.frontlineonnet.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'traveller.outlookindia.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'www.thehindu.com', 'books.google.com', 'timesofindia.indiatimes.com', 'timesmachine.nytimes.com', 'books.google.com', 'www.youtube.com', 'www.cookawesome.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.youtube.com', 'books.google.com', 'books.google.com', 'english.manoramaonline.com', 'www.thetakeiteasychef.com', 'books.google.com', 'www.facesplacesandplates.com', 'www.frontlineonnet.com', 'www.outlookindia.com', 'books.google.com', 'www.hindu.com', 'books.google.com', 'books.google.com', 'www.kozhikodeairport.com', 'books.google.com', 'www.gutenberg.org', 'worldcat.org', ['muallim journal of social sciences and humanities']]",1574251,Allow all users (no expiry set),68478,6 March 2005,QuartierLatin1968 ,1399,10,2005-03-06,2005-03,2005
484,484,Culture of the Song dynasty,https://en.wikipedia.org/wiki/Culture_of_the_Song_dynasty,90,0,[],[],0,0,0,1,0,0,89,0.0,0.0,0.011111111111111112,0.0,0.0,0.0,0,['arts.cultural-china.com'],10443917,Allow all users (no expiry set),72197,3 April 2007,PericlesofAthens ,698,0,2007-04-03,2007-04,2007
485,485,Arbëreshë people,https://en.wikipedia.org/wiki/Arb%C3%ABresh%C3%AB_people,31,2,"['10.1038/s41598-017-01802-4', '10.1515/ijsl.2006.014', '28512355', None, '5434004', None]","[['scientific reports '], [' international journal of the sociology of language']]",1,0,0,14,0,0,14,0.03225806451612903,0.0,0.45161290322580644,0.06451612903225806,0.0,0.0967741935483871,2,"['search.proquest.com', 'books.google.com', 'lulu.com', 'search.proquest.com', 'www.ethnologue.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.nature.com', 'www.insajderi.com', 'benjamins.com', 'books.google.com', 'books.google.com', 'lucania1.altervista.org', ['scientific reports '], [' international journal of the sociology of language']]",429498,Allow all users (no expiry set),46294,13 January 2004,213.103.134.167 ,1458,2,2004-01-13,2004-01,2004
486,486,Rajbiraj,https://en.wikipedia.org/wiki/Rajbiraj,74,0,[],[],3,6,0,51,0,0,14,0.04054054054054054,0.08108108108108109,0.6891891891891891,0.0,0.0,0.12162162162162163,0,"['www.rajbirajmun.gov', 'www.dhm.gov', 'cbs.gov', 'www.rajbirajmun.gov', 'cbs.gov', 'www.moic.gov', 'bossnepal.com', 'rajbirajdainik.com', 'books.google.com', 'www.onlinekhabar.com', 'www.goalnepal.com', 'nagariknews.nagariknetwork.com', 'thehimalayantimes.com', 'thehimalayantimes.com', 'www.myrepublica.com', 'deshsanchar.com', 'www.republicadainik.com', 'cricketingnepal.com', 'myrepublica.nagariknetwork.com', 'thehimalayantimes.com', 'archive.nepalitimes.com', 'www.spotlightnepal.com', 'books.google.com', 'myrepublica.nagariknetwork.com', 'kathmandupost.com', 'trn.gorkhapatraonline.com', 'myrepublica.nagariknetwork.com', 'google.com', 'www.sites.google.com', 'thehimalayantimes.com', 'thehimalayantimes.com', 'www.collegenp.com', 'myrepublica.nagariknetwork.com', 'www.asianart.com', 'ekantipur.com', 'newstoday.com', 'www.hakahaki.com', 'www.buddhaair.com', 'myrepublica.com', 'books.google.com', 'nepalitimes.com', 'kathmandupost.com', 'www.housingnepal.com', 'newstoday.com', 'myrepublica.nagariknetwork.com', 'kathmandupost.com', 'ekantipur.com', 'kathmandupost.ekantipur.com', 'kathmandupost.ekantipur.com', 'kathmandupost.com', 'newstoday.com', 'www.majheri.com', 'thehimalayantimes.com', 'thehimalayantimes.com', 'www.spotlightnepal.com', 'kathmandupost.com', 'thehimalayantimes.com', 'www.madanpuraskar.org', 'unstats.un.org', 'www.therisingnepal.org']",1270030,Allow all users (no expiry set),41613,12 December 2004,217.43.194.58 ,711,0,2004-12-12,2004-12,2004
487,487,Southern Serbia (geographical region),https://en.wikipedia.org/wiki/Southern_Serbia_(geographical_region),24,0,[],[],4,2,0,5,0,0,13,0.16666666666666666,0.08333333333333333,0.20833333333333334,0.0,0.0,0.25,0,"['stat.gov', 'crm.siepa.gov', 'kraljevo-cafe.com', 'www.juznevesti.com', 'www.juznevesti.com', 'sacred-texts.com', 'www.juznevesti.com', 'unesco.org', 'www.centenaire.org', 'unesco.org', 'www.makroekonomija.org']",66169508,Allow all users (no expiry set),28154,21 December 2020,SRofSerbia ,58,1,2020-12-21,2020-12,2020
488,488,List of English words of French origin,https://en.wikipedia.org/wiki/List_of_English_words_of_French_origin,3,0,[],[],0,0,0,2,0,0,1,0.0,0.0,0.6666666666666666,0.0,0.0,0.0,0,"['www.connexionfrance.com', 'www.connexionfrance.com']",566269,Allow all users (no expiry set),29119,31 March 2004,Fabiform ,1765,2,2004-03-31,2004-03,2004
489,489,Newar people,https://en.wikipedia.org/wiki/Newar_people,129,2,"['10.24924/ijise/2017.04/v5.iss2/1.12', '10.2307/2843991', None, None, None, None]","[['international journal of information systems and engineering'], [' journal of the royal anthropological institute', 'royal anthropological institute of great britain and ireland']]",19,6,0,44,0,1,57,0.14728682170542637,0.046511627906976744,0.34108527131782945,0.015503875968992248,0.0,0.20930232558139536,2,"['cbs.gov', 'www.kathmandu.gov', 'cbs.gov', 'www.cbs.gov', 'www.cbs.gov', 'cbs.gov', 'web.com', 'nationalgeographic.com', 'web.com', 'www.ekantipur.com', 'www.thehimalayantimes.com', 'www.nepalitimes.com', 'cis.sagepub.com', 'newaissues.wordpress.com', 'www.sothebys.com', 'web.com', 'www.kpmalla.com', 'www.dancemandal.com', 'web.com', 'www.kpmalla.com', 'books.google.com', 'www.digitalhimalaya.com', 'books.google.com', 'dictionary.reference.com', 'books.google.com', 'e.myrepublica.com', 'thehimalayantimes.com', 'www.kpmalla.com', 'www.kpmalla.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'thehimalayantimes.com', 'cis.sagepub.com', 'books.google.com', 'www.kpmalla.com', 'books.google.com', 'web.com', 'e.myrepublica.com', 'www.kpmalla.com', 'www.scribd.com', 'buddhim.20m.com', 'www.facebook.com', 'www.artsofnepal.com', 'www.kpmalla.com', 'www.digitalhimalaya.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'www.kpmalla.com', 'seechac.org', 'unesdoc.unesco.org', 'publishing.cdlib.org', 'www.gutenberg.org', 'journals.cambridge.org', 'publishing.cdlib.org', 'unesdoc.unesco.org', 'www.newarsinsikkim.org', 'www.ppguk.org', 'www.gutenberg.org', 'www.gutenberg.org', 'www.anuttaratrikakula.org', 'www.gutenberg.org', 'unesdoc.unesco.org', 'unesdoc.unesco.org', 'www.newajapan.org', 'whc.unesco.org', 'www.newah.org', 'www.gutenberg.org', ['international journal of information systems and engineering'], [' journal of the royal anthropological institute', 'royal anthropological institute of great britain and ireland']]",997963,Allow all users (no expiry set),80406,19 September 2004,Alberuni ,1533,11,2004-09-19,2004-09,2004
490,490,Kashubians,https://en.wikipedia.org/wiki/Kashubians,70,5,"['10.1371/journal.pone.0054360', '10.1038/ejhg.2012.190', '10.1080/00905999708408536', '10.1371/journal.pone.0135820', '10.1002/ajpa.21253', '23342138', '22968131', None, '26332464', '20091807', '3544712', '3598329', None, '4558026', None]","[['[[plos one'], ['european journal of human genetics'], [' [[nationalities papers'], ['[[plos one'], ['[[american journal of physical anthropology']]",3,5,0,6,0,0,51,0.04285714285714286,0.07142857142857142,0.08571428571428572,0.07142857142857142,0.0,0.18571428571428572,5,"['www.stat.gov', 'www.senat.gov', 'www.gov', 'stat.gov', 'www.stat.gov', 'findarticles.com', 'kaszebsko.com', 'www.worldatlas.com', 'www.omniglot.com', 'books.google.com', 'kaszebsko.com', 'bambenek.org', 'uu.diva-portal.org', 'bambenek.org', ['[[plos one'], ['european journal of human genetics'], [' [[nationalities papers'], ['[[plos one'], ['[[american journal of physical anthropology']]",17020,Allow all users (no expiry set),57240,17 October 2001,Rmhermen ,1108,1,2001-10-17,2001-10,2001
491,491,Jianghuai people,https://en.wikipedia.org/wiki/Jianghuai_people,16,0,[],[],0,0,0,7,0,0,9,0.0,0.0,0.4375,0.0,0.0,0.0,0,"['www.chinatouradvisors.com', 'www.statista.com', 'www.zhonghuashu.com', 'www.zhonghuashu.com', 'www.ziyexing.com', 'www.theworldofchinese.com', 'sfrichmondreview.com']",54636085,Allow all users (no expiry set),17354,24 July 2017,Kamikaze2017 ,129,1,2017-07-24,2017-07,2017
492,492,Larissa,https://en.wikipedia.org/wiki/Larissa,32,0,[],[],2,2,0,1,0,0,27,0.0625,0.0625,0.03125,0.0,0.0,0.125,0,"['www.larissa.gov', 'ftp.atdd.noaa.gov', 'www.larissa.climatemps.com', 'plato-dialogues.org', 'meteo-climat-bzh.dyndns.org']",18490,Allow all users (no expiry set),45616,30 November 2001,Bryan Derksen ,1634,2,2001-11-30,2001-11,2001
493,493,Gujarati people,https://en.wikipedia.org/wiki/Gujarati_people,215,5,"['10.1080/14736489.2016.1165557', '10.2307/1166488', '10.1057/9781403914484_4', '10.3765/bls.v36i1.3917', '10.2307/2060606', None, None, None, None, '5163987', None, None, None, None, None]","[['[[taylor ', 'india review'], ['issue'], ['palgrave macmillan'], ['annual meeting of the berkeley linguistics society'], ['demography']]",11,6,0,154,0,0,39,0.05116279069767442,0.027906976744186046,0.7162790697674418,0.023255813953488372,0.0,0.10232558139534884,5,"['www.dhs.gov', 'www.dhs.gov', 'www.dhs.gov', 'www.dhs.gov', 'uidai.gov', 'www.stats.gov', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'www.thenews.com', 'alivelshi.com', 'bollyspice.com', 'blogs.timesofindia.indiatimes.com', 'www.nytimes.com', 'www.newindianexpress.com', 'books.google.com', 'www.jaincentreleicester.com', 'www.nybooks.com', 'books.google.com', 'books.google.com', 'nonconformer.wordpress.com', 'www.perthnow.com', 'mangalayatan.com', 'mayamovies.com', 'timesofindia.indiatimes.com', 'www.facebook.com', 'www.economist.com', 'books.google.com', 'www.torontogarba.com', 'timesofindia.indiatimes.com', 'articles.economictimes.indiatimes.com', 'photogallery.indiatimes.com', 'books.google.com', 'www.magepublishers.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.rogerebert.com', 'timesofindia.indiatimes.com', 'www.rhcapitalpartners.com', 'books.google.com', 'timesofindia.indiatimes.com', 'espncricinfo.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'sklpc.com', 'books.google.com', 'profile.id.com', 'articles.economictimes.indiatimes.com', 'books.google.com', 'dnaindia.com', 'www.td.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.businessdailyafrica.com', 'www.thehindu.com', 'books.google.com', 'theconversation.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'm.timesofindia.com', 'www.facebook.com', 'www.gujaratimuslimmarriage.com', 'books.google.com', 'books.google.com', 'india.blogs.nytimes.com', 'cineplot.com', 'deshgujarat.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.td.com', 'timesofindia.indiatimes.com', 'blogs.wsj.com', 'timesofindia.indiatimes.com', 'www.thestar.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'zeenews.india.com', 'parthoza.com', 'timesofindia.indiatimes.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.facebook.com', 'books.google.com', 'www.facebook.com', 'books.google.com', 'books.google.com', 'books.google.com', 'theindiandiaspora.com', 'www.khanakhazana.com', 'www.karismatickarachi.com', 'timesofindia.indiatimes.com', 'www.bhatiamahajan.com', 'business.in.com', 'www.bollywoodlife.com', 'books.google.com', 'timesofindia.indiatimes.com', 'pressreader.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'www.businessdailyafrica.com', 'timesofindia.indiatimes.com', 'www.canada.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thenews.com', 'timesofindia.indiatimes.com', 'alusainc.wordpress.com', 'timesofindia.indiatimes.com', 'www.bloomberg.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'thestar.com', 'books.google.com', 'blogs.economictimes.indiatimes.com', 'tribune.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.sfgate.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thenews.com', 'books.google.com', 'books.google.com', 'www.indiaglitz.com', 'buddybits.com', 'deshgujarat.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.kenyanentrepreneur.com', 'books.google.com', 'www.intlgymnast.com', 'articles.economictimes.indiatimes.com', 'timesofindia.indiatimes.com', 'books.google.com', 'outlookindia.com', 'www.dnaindia.com', 'rediff.com', 'books.google.com', 'books.google.com', 'nymag.com', 'books.google.com', 'books.google.com', 'blog.mapsofindia.com', 'ndtv.com', 'timesofindia.indiatimes.com', 'www.sahistory.org', 'sahistory.org', 'sahistory.org', 'www.rajsaubhag.org', 'natalia.org', 'www.countercurrents.org', 'www.jstor.org', 'maheronline.org', 'www.natalia.org', 'ukncgo.org', 'www.eauk.org', ['[[taylor ', 'india review'], ['issue'], ['palgrave macmillan'], ['annual meeting of the berkeley linguistics society'], ['demography']]",6320523,Allow all users (no expiry set),145955,20 July 2005,BD2412 ,4210,52,2005-07-20,2005-07,2005
494,494,Culture of the Czech Republic,https://en.wikipedia.org/wiki/Culture_of_the_Czech_Republic,16,1,"['10.1387/veleia.18074', None, None]",[['veleia ']],4,0,0,4,0,0,7,0.25,0.0,0.25,0.0625,0.0,0.3125,1,"['www.archdaily.com', 'www.nytimes.com', 'worldpopulationreview.com', 'www.bbc.com', 'nobelprize.org', 'whc.unesco.org', 'awardsdatabase.oscars.org', 'nobelprize.org', ['veleia ']]",6675817,Allow all users (no expiry set),15825,25 August 2006,Jax-wp ,272,0,2006-08-25,2006-08,2006
495,495,Syrians,https://en.wikipedia.org/wiki/Syrians,125,12,"['10.1086/511103', '10.1126/science.290.5494.1155', '10.1371/journal.pone.0054616', '10.1073/pnas.100115997', '10.1111/j.1469-1809.2009.00538.x', '10.1086/373570', '10.1038/srep35837', '10.1371/journal.pgen.1003316', '10.1371/journal.pone.0118625', '10.1038/ejhg.2010.177', '10.3406/topoi.2009.2306', '10.1371/journal.pone.0192269', None, '11073453', '23382925', '10801975', '19686289', None, '27848937', '23468648', '25738654', '21119711', None, '29522542', None, None, '3559847', '18733', '3312577', None, '5111078', '3585000', '4349752', '3062011', None, '5844529']","[['journal of near eastern studies '], ['science '], ['plos one'], ['pnas', ' proceedings of the national academy of sciences'], [' annals of human genetics'], ['journal of near eastern studies '], ['scientific reports '], [' plos genetics '], ['plos one'], ['european journal of human genetics'], ['topoi. orient-occident', 'société des amis de la bibliothèque salomon-reinach'], ['plos one']]",11,5,0,33,0,0,64,0.088,0.04,0.264,0.096,0.0,0.224,12,"['factfinder.census.gov', 'cia.gov', 'www.itamaraty.gov', 'state.gov', 'www.cia.gov', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.businessweek.com', 'books.google.com', 'books.google.com', 'caribbeanhistoryarchives.blogspot.com', 'www.forbes.com', 'arabnews.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.newyorker.com', 'books.google.com', 'jusoorsyria.com', 'www.thaindian.com', 'books.google.com', 'books.google.com', 'aawsat.com', 'www.bloomberg.com', 'www.wamda.com', 'www.forbes.com', 'books.google.com', 'priyadsouza.com', 'gulfnews.com', 'books.google.com', 'www.businessweek.com', 'books.google.com', 'iberoamericasocial.com', 'books.google.com', 'www.reuters.com', 'pomeps.org', 'unhcr.org', 'data2.unhcr.org', 'unhcr.org', 'www.jaas.org', 'www.as-coa.org', 'www.ieee-ras.org', 'aristobulo.psuv.org', 'data2.unhcr.org', 'unhcr.org', 'amerika.revues.org', ['journal of near eastern studies '], ['science '], ['plos one'], ['pnas', ' proceedings of the national academy of sciences'], [' annals of human genetics'], ['journal of near eastern studies '], ['scientific reports '], [' plos genetics '], ['plos one'], ['european journal of human genetics'], ['topoi. orient-occident', 'société des amis de la bibliothèque salomon-reinach'], ['plos one']]",8862873,Allow all users (no expiry set),79565,11 January 2007,Beland ,1735,13,2007-01-11,2007-01,2007
496,496,Faisalabad,https://en.wikipedia.org/wiki/Faisalabad,190,1,"['10.1073/pnas.1112743109', '22645375', '3387054']","[['pnas', 'national academy of sciences ']]",17,40,0,88,0,0,44,0.08947368421052632,0.21052631578947367,0.4631578947368421,0.005263157894736842,0.0,0.30526315789473685,1,"['www.urbanunit.gov', 'faisalabad.gov', 'www.radio.gov', 'www.faisalabad.gov', 'punjab.gov', 'fwf.punjab.gov', 'faisalabad.gov', 'namc.pmd.gov', 'www.railways.gov', 'www.faisalabadpolice.gov', 'www.pmd.gov', 'www.pta.gov', 'punjab.gov', 'prr.hec.gov', 'www.dgtrdt.gov', 'www.fwf.punjab.gov', 'faisalabadpolice.gov', 'pbs.gov', 'www.faisalabad.gov', 'www.punjab.gov', 'www.pmd.gov', 'rmcpunjab.pmd.gov', 'prr.hec.gov', 'faisalabad.dc.lhc.gov', 'www.hec.gov', 'www.pemra.gov', 'namc.pmd.gov', 'www.cm.punjab.gov', 'nha.gov', 'www.pta.gov', 'faisalabad.dc.lhc.gov', 'faisalabad.dc.lhc.gov', 'www.faisalabadartscouncil.gov', 'www.punjab.gov', 'www.radio.gov', 'punjablaws.gov', 'lgcd.punjab.gov', 'www.punjab.gov', 'faisalabad.gov', 'fwf.punjab.gov', 'www.pakistantoday.com', 'www.thenews.com', 'nation.com', 'fiedmc.com', 'tribune.com', 'www.serenahotels.com', 'nation.com', 'www.dawn.com', 'www.dawn.com', 'tribune.com', 'tribune.com', 'tribune.com', 'www.bbc.com', 'www.pakladies.com', 'tribune.com', 'books.google.com', 'www.embassypages.com', 'tribune.com', 'www.gulfair.com', 'books.google.com', 'www.caapakistan.com', 'tribune.com', 'books.google.com', 'www.foxnews.com', 'www.highbeam.com', 'www.thenews.com', 'books.google.com', 'www.urdupoint.com', 'www.washingtonpost.com', 'tribune.com', 'books.google.com', 'pakistaniat.com', 'books.google.com', 'www.asian-recipe.com', 'books.google.com', 'cricketarchive.com', 'www.pakistanitourism.com', 'ndtvsports.com', 'www.britannica.com', 'www.thenewstribe.com', 'www.urdupoint.com', 'www.subrung.com', 'www.youtube.com', 'fcci.com', 'tribune.com', 'www.dailytimes.com', 'tribune.com', 'chenabclub.com', 'www.fcci.com', 'tribune.com', 'www.brecorder.com', 'books.google.com', 'citypulse.com', 'tribune.com', 'tribune.com', 'www.atimes.com', 'www.thenews.com', 'tribune.com', 'www.dawn.com', 'www.scribd.com', 'books.google.com', 'www.lawsofpakistan.com', 'www.pakimag.com', 'ptcl.com', 'www.pakmet.com', 'dawn.com', 'www.fcci.com', 'nation.com', 'tribune.com', 'cinenagina.com', 'www.fcci.com', 'tribune.com', 'nation.com', 'books.google.com', 'www.cinepax.com', 'www.qatarairways.com', 'www.dawn.com', 'cricketarchive.com', 'www.nespak.com', 'www.espncricinfo.com', 'faisalabad.com', 'www.thenews.com', 'tribune.com', 'www.bloomberg.com', 'www.journeum.com', 'nation.com', 'books.google.com', 'www.youtube.com', 'www.npr.org', 'www.pakistanpressfoundation.org', 'www.jstor.org', 'www.ijser.org', 'www.asb.org', 'pwon.org', 'www.smeda.org', 'www.aserpakistan.org', 'www.wto.org', 'agris.fao.org', 'www.internews.org', 'faisalabadliteraryfestival.org', 'www.asb.org', 'unesco.org', 'pakvoter.org', 'climate-data.org', 'www.flaginstitute.org', ['pnas', 'national academy of sciences ']]",401880,Allow all users (no expiry set),111163,14 December 2003,ThaGrind ,5295,14,2003-12-14,2003-12,2003
497,497,Nafplio,https://en.wikipedia.org/wiki/Nafplio,38,0,[],[],0,0,0,6,0,0,32,0.0,0.0,0.15789473684210525,0.0,0.0,0.0,0,"['books.google.com', 'visitnafplio.com', 'query.nytimes.com', 'ypodomes.com', 'www.menton.com', 'www.vniles.com']",966904,Allow all users (no expiry set),30478,7 September 2004,Mozzerati ,557,0,2004-09-07,2004-09,2004
498,498,Christian culture,https://en.wikipedia.org/wiki/Christian_culture,346,12,"['10.2307/1291170', None, '10.1057/9781403980618', '10.1017/cbo9780511676062', '10.1080/08873630802617135', '10.2307/1952449', '10.1353/jhi.2006.0035', '10.1080/10253860500160361', '10.1093/acref/9780198607663.001.0001', '10.1111/j.1467-9558.2009.01367.x', '10.1162/0022195052564243', '10.1080/14650040903420388', None, '3902734', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None]","[['dumbarton oaks papers', 'dumbarton oaks'], ['the henry e. sigerist supplements to the bulletin of the history of medicine', 'johns hopkins'], ['palgrave macmillan '], [' cambridge university press '], ['journal of cultural geography', ' routledge'], ['[[american political science review'], ['journal of the history of ideas '], ['consumption markets '], ['oxford university press '], [' sociological theory '], [' the journal of interdisciplinary history'], ['geopolitics']]",29,2,0,94,0,3,207,0.0838150289017341,0.005780346820809248,0.27167630057803466,0.03468208092485549,0.0,0.12427745664739884,12,"['www.opm.gov', 'www.direct.gov', 'www.adherents.com', 'content.time.com', 'www.eotc.faithweb.com', 'books.google.com', 'www.guinnessworldrecords.com', 'www.christiansofiraq.com', 'www.vanityfair.com', 'www.nytimes.com', 'books.google.com', 'www.sfgate.com', 'www.german-way.com', 'books.google.com', 'books.google.com', 'books.google.com', 'boxofficemojo.com', 'www.touchstonemag.com', 'diepresse.com', 'www.britannica.com', 'en.biginfinland.com', 'search.ebscohost.com', 'books.google.com', 'books.google.com', 'www.washingtonpost.com', 'books.google.com', 'www.britannica.com', 'www.britannica.com', 'miradaglobal.com', 'about.com', 'www.britannica.com', 'www.siouxcityjournal.com', 'books.google.com', 'www.infoplease.com', 'www.gallup.com', 'books.google.com', 'www.dictionaryofchristianese.com', 'issuu.com', 'www.nbcnews.com', 'www.nbcnews.com', 'books.google.com', 'books.google.com', 'www.touchstonemag.com', 'books.google.com', 'insidemovies.moviefone.com', 'www.catholicnewsagency.com', 'historymedren.about.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.creationsafaris.com', 'www.adherents.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.boxofficemojo.com', 'www.nrbookservice.com', 'books.google.com', 'www.economist.com', 'books.google.com', 'variety.com', 'www.britannica.com', 'www.adherents.com', 'www.deseretnews.com', 'books.google.com', 'www.goodreads.com', 'www.britannica.com', 'books.google.com', 'www.ewtn.com', 'www.onlinedigeditions.com', 'nippon.com', 'books.google.com', 'college.hmco.com', 'books.google.com', 'www.britannica.com', 'www.britannica.com', 'www.deseretnews.com', 'adherents.com', 'books.google.com', 'www.nytimes.com', 'www.boxofficemojo.com', 'books.google.com', 'www.christianpost.com', 'timesmachine.nytimes.com', 'www.time.com', 'books.google.com', 'www.turkmenhost.com', 'books.google.com', 'books.google.com', 'www.ewtn.com', 'books.google.com', 'www.britannica.com', 'www.wsj.com', 'www.adherents.com', 'www.adherents.com', 'adherents.com', 'www.pewforum.org', 'www.newadvent.org', 'www.godandscience.org', 'www.chesterton.org', 'religion-online.org', 'www.malayalamresourcecentre.org', 'www.salvationarmy-newyork.org', 'pnclink.org', 'www.chesterton.org', 'biologos.org', 'www.middle-ages.org', 'assets.pewresearch.org', 'www.pewforum.org', 'www.worldcat.org', 'www.newadvent.org', 'newadvent.org', 'newadvent.org', 'broughttolife.sciencemuseum.org', 'archives.umc.org', 'newadvent.org', 'www.pewresearch.org', 'www.doaks.org', 'www.usccb.org', 'www.pewforum.org', 'www.churchofjesuschrist.org', 'rae.org', 'openlibrary.org', 'www.catholiceducation.org', 'www.newadvent.org', ['dumbarton oaks papers', 'dumbarton oaks'], ['the henry e. sigerist supplements to the bulletin of the history of medicine', 'johns hopkins'], ['palgrave macmillan '], [' cambridge university press '], ['journal of cultural geography', ' routledge'], ['[[american political science review'], ['journal of the history of ideas '], ['consumption markets '], ['oxford university press '], [' sociological theory '], [' the journal of interdisciplinary history'], ['geopolitics']]",32516987,Allow all users (no expiry set),216056,24 July 2011,Dbachmann ,366,2,2011-07-24,2011-07,2011
499,499,Pontremoli,https://en.wikipedia.org/wiki/Pontremoli,13,0,[],[],0,0,0,9,0,1,3,0.0,0.0,0.6923076923076923,0.0,0.0,0.0,0,"['www.britannica.com', 'www.com', 'books.google.com', 'www.wsj.com', 'books.google.com', 'about.com', 'www.wsj.com', 'www.britannica.com', 'books.google.com']",4067694,Allow all users (no expiry set),13084,14 February 2006,Bogdangiusca ,205,1,2006-02-14,2006-02,2006
500,500,Galilee,https://en.wikipedia.org/wiki/Galilee,29,0,[],[],4,3,0,13,0,0,9,0.13793103448275862,0.10344827586206896,0.4482758620689655,0.0,0.0,0.2413793103448276,0,"['www.cbs.gov', 'www.cbs.gov', 'www.cbs.gov', 'ancienthistory.about.com', 'www.govisitisrael.com', 'books.google.com', 'ca.news.yahoo.com', 'www.jewishsf.com', 'books.google.com', 'sciencedaily.com', 'books.google.com', 'books.google.com', 'ynetnews.com', 'books.google.com', 'fr.jpost.com', 'www.dictionary.com', 'data.perseus.org', 'www.jafi.org', 'www.jta.org', 'jewishvirtuallibrary.org']",12639,Require extended confirmed access (no expiry set),38997,29 September 2001,216.99.203.xxx ,1088,0,2001-09-29,2001-09,2001
501,501,Coimbatore district,https://en.wikipedia.org/wiki/Coimbatore_district,109,1,"['10.11609/jott.zpj.1657.2944-8', None, None]",[['zoos']],2,9,0,80,0,0,17,0.01834862385321101,0.08256880733944955,0.7339449541284404,0.009174311926605505,0.0,0.11009174311926606,1,"['www.tn.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'www.ccmc.gov', 'www.tn.gov', 'www.censusindia.gov', 'pibmumbai.gov', 'www.censusindia.gov', 'www.tn.gov', 'books.google.com', 'hindu.com', 'www.hinduonnet.com', 'www.thehindubusinessline.com', 'www.hindustantimes.com', 'www.deccanchronicle.com', 'articles.timesofindia.indiatimes.com', 'www.thehindubusinessline.com', 'www.hindu.com', 'www.hinduonnet.com', 'www.hindu.com', 'www.thecityvisit.com', 'www.hindu.com', 'www.hindu.com', 'www.resourceinvestor.com', 'www.hindu.com', 'www.hinduonnet.com', 'www.resourceinvestor.com', 'www.hinduonnet.com', 'siliconindia.com', 'articles.timesofindia.indiatimes.com', 'www.thehindu.com', 'www.hinduonnet.com', 'www.thehindubusinessline.com', 'www.ndtv.com', 'www.thehindubusinessline.com', 'www.hindu.com', 'articles.economictimes.indiatimes.com', 'tamil.dinamalar.com', 'www.thehindu.com', 'mydigitalfc.com', 'www.hindu.com', 'www.exchange4media.com', 'smetimes.tradeindia.com', 'www.thehindubusinessline.com', 'archive.financialexpress.com', 'articles.timesofindia.indiatimes.com', 'thehindujobs.com', 'indiaprwire.com', 'www.vivantabytaj.com', 'books.google.com', 'www.hindu.com', 'books.google.com', 'commodityonline.com', 'news.google.com', 'www.winentrance.com', 'www.hindu.com', 'www.hindu.com', 'economictimes.indiatimes.com', 'www.hindu.com', 'www.hinduonnet.com', 'www.thehindu.com', 'www.thehindu.com', 'www.hinduonnet.com', 'www.hindu.com', 'www.hindu.com', 'www.hindu.com', 'www.moneycontrol.com', 'intecexpo.com', 'www.hindu.com', 'www.hindu.com', 'o3.indiatimes.com', 'www.thehindu.com', 'www.hindu.com', 'newindianexpress.com', 'www.hindu.com', 'timesofindia.indiatimes.com', 'www.moneycontrol.com', 'timesofindia.indiatimes.com', 'eproceedings.worldscinet.com', 'www.hindu.com', 'www.hindu.com', 'www.hindu.com', 'www.hindu.com', 'www.hinduonnet.com', 'tamilnadu.com', 'www.thehindu.com', 'www.thehindubusinessline.com', 'www.thehindu.com', 'www.thehindu.com', 'govartcbe.org', 'whc.unesco.org', ['zoos']]",3829700,Allow all users (no expiry set),74136,24 January 2006,Cheeni ,960,4,2006-01-24,2006-01,2006
502,502,Pathans in India,https://en.wikipedia.org/wiki/Pathans_in_India,157,0,[],[],7,2,0,135,0,0,13,0.044585987261146494,0.012738853503184714,0.8598726114649682,0.0,0.0,0.05732484076433121,0,"['prasarbharati.gov', 'censusindia.gov', 'livemint.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.ndtv.com', 'www.aljazeera.com', 'www.business-standard.com', 'www.youtube.com', 'books.google.com', 'www.rediff.com', 'books.google.com', 'books.google.com', 'dailytimes.com', 'tribune.com', 'books.google.com', 'tribune.com', 'books.google.com', 'books.google.com', 'www.hindustantimes.com', 'www.dawn.com', 'www.dawn.com', 'www.seattlepi.com', 'indianexpress.com', 'books.google.com', 'www.outlookindia.com', 'muslimmirror.com', 'books.google.com', 'www.nytimes.com', 'www.wionews.com', 'books.google.com', 'www.rediff.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'www.tribuneindia.com', 'www.sentinelassam.com', 'tribune.com', 'books.google.com', 'books.google.com', 'www.outlookindia.com', 'newsonair.com', 'books.google.com', 'www.thesundayindian.com', 'books.google.com', 'books.google.com', 'dailytimes.com', 'books.google.com', 'www.cinestaan.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.outlookindia.com', 'books.google.com', 'www.britannica.com', 'www.thehindu.com', 'www.thehindu.com', 'www.deccanherald.com', 'indianexpress.com', 'www.hindustantimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.bbc.com', 'food.ndtv.com', 'www.dawn.com', 'www.newindianexpress.com', 'books.google.com', 'www.thehindubusinessline.com', 'www.youtube.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thebetterindia.com', 'www.deccanherald.com', 'www.newindianexpress.com', 'books.google.com', 'openthemagazine.com', 'books.google.com', 'photogallery.indiatimes.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'www.thenews.com', 'books.google.com', 'www.hindustantimes.com', 'books.google.com', 'books.google.com', 'qz.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'www.aljazeera.com', 'zeenews.india.com', 'books.google.com', 'books.google.com', 'www.dnaindia.com', 'www.business-standard.com', 'food.ndtv.com', 'www.thecrimson.com', 'openthemagazine.com', 'www.hindustantimes.com', 'books.google.com', 'www.rediff.com', 'books.google.com', 'www.hindustantimes.com', 'www.dailytimes.com', 'www.hindustantimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'indianexpress.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'www.ussquash.com', 'books.google.com', 'www.hindustantimes.com', 'www.tribuneindia.com', 'www.hindustantimes.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'punemirror.indiatimes.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.thenews.com', 'indianexpress.com', 'www.dawn.com', 'books.google.com', 'khyber.org', 'en.banglapedia.org', 'www.bharatiyahockey.org', 'guyana.org', 'www.afghanistan-analysts.org', 'www.jstor.org', 'airworldservice.org']",64100474,Allow all users (no expiry set),95592,28 May 2020,Mar4d ,466,7,2020-05-28,2020-05,2020
503,503,Andalusia,https://en.wikipedia.org/wiki/Andalusia,213,4,"['10.1163/157006709x458891', '10.1515/islm.1989.66.2.252', '10.12795/rea.1986.i07.02', '10.1086/467294', None, None, None, None, None, None, None, None]","[['medieval encounters', 'brill nv'], ['der islam'], [' revista de estudios andaluces'], ['[[the journal of law and economics']]",11,1,0,43,0,0,154,0.051643192488262914,0.004694835680751174,0.20187793427230047,0.018779342723004695,0.0,0.07511737089201878,4,"['estatico.buenosaires.gov', 'books.google.com', 'www.antonioburgos.com', 'www.lavanguardia.com', 'renewableenergymagazine.com', 'www.flamenco-world.com', 'books.google.com', 'books.google.com', 'books.google.com', 'hermandadrociosevilla.com', 'www.elpais.com', 'www.energias-renovables.com', 'www.andaluciafilm.com', 'books.google.com', 'fórmulatv.com', 'andalucia.com', 'www.andaluciainvestiga.com', 'abodeinternational.com', 'www.collinsdictionary.com', 'visithuelva.com', 'www.mocavo.com', 'cervantesvirtual.com', 'en.oxforddictionaries.com', 'books.google.com', 'www.myhomeinandalucia.com', 'www.andalucia.com', 'files.shareholder.com', 'www.valemusic.com', 'uefa.com', 'www.myhomeinandalucia.com', 'www.iberianature.com', 'books.google.com', 'www.iberianature.com', 'www.andalucia.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.jotamartin.byethost33.com', 'noticias.juridicas.com', 'books.google.com', 'ecoticias.com', 'books.google.com', 'www.correodelmaestro.com', 'www.britannica.com', 'www.accessibletourism.org', 'es.wikisource.org', 'archnet.org', 'www.fundacionandaluciaolimpica.org', 'es.climate-data.org', 'www.andalucia.org', 'www.ecologistasenaccion.org', 'www.fttcv.org', 'www.fao.org', 'www.realescuela.org', 'sustainabletourismworld.org', ['medieval encounters', 'brill nv'], ['der islam'], [' revista de estudios andaluces'], ['[[the journal of law and economics']]",2736,Allow all users (no expiry set),218506,29 November 2001,Tsja ,3289,6,2001-11-29,2001-11,2001
504,504,Međimurje County,https://en.wikipedia.org/wiki/Me%C4%91imurje_County,12,0,[],[],1,0,0,1,0,0,10,0.08333333333333333,0.0,0.08333333333333333,0.0,0.0,0.08333333333333333,0,"['www.mtraditional.com', 'hdi.globaldatalab.org']",435781,Allow all users (no expiry set),50174,19 January 2004,68.249.230.114 ,1478,0,2004-01-19,2004-01,2004
505,505,Islam in Uttar Pradesh,https://en.wikipedia.org/wiki/Islam_in_Uttar_Pradesh,43,0,[],[],2,1,0,11,0,0,29,0.046511627906976744,0.023255813953488372,0.2558139534883721,0.0,0.0,0.06976744186046512,0,"['www.censusindia.gov', 'www.deccanherald.com', 'szh.20m.com', 'www.geocities.com', 'www.britannica.com', 'www.questia.com', 'articles.timesofindia.indiatimes.com', 'books.google.com', 'www.languageinindia.com', 'theurdulanguage.com', 'india_resource.tripod.com', 'india_resource.tripod.com', 'www.ethnologue.org', 'muslimsocieties.org']",28257071,Allow all users (no expiry set),44895,4 August 2010,WALTHAM2 ,515,2,2010-08-04,2010-08,2010
506,506,List of Italian inventions and discoveries,https://en.wikipedia.org/wiki/List_of_Italian_inventions_and_discoveries,571,57,"['10.1111/j.1600-0773.1948.tb03345.x', '10.5951/mt.57.5.0323', '10.1056/nejmp030080', '10.1038/nature.2017.22231', '10.1002/clc.4960251010', '10.1109/mpe.2007.904752', '10.1038/280707a0', '10.1051/epjconf/201714302149', '10.4000/archeomed.18586', '10.1016/j.nlm.2017.04.010', '10.2307/3100858', '10.1007/bf01696201', '10.1038/366716b0', '10.5152/balkanmedj.2013.003', '10.1073/pnas.1324149111', '10.1097/01.brs.0000182314.49515.d8', '10.5642/perfpr.201318.01.05', '10.1016/s0893-133x(99)00031-7', None, '10.1016/s0141-3910(97)00156-0', '10.3762/bjnano.4.37', None, '10.2307/3574319', '10.1172/jci77540', '10.1177/003591573002300445', '10.1227/01.neu.0000139458.36781.31', '10.1080/10623320802092377', '10.1103/physrev.54.772.2', '10.1016/s0262-4079(10)62415-3', '10.1084/jem.20151960', '10.1097/00007632-200001010-00022', '10.1103/physrev.58.672', '10.1103/physreva.65.062710', '10.2307/4344123', None, '10.1016/s0065-2164(01)48005-1', '10.1038/159024a0', '10.1103/physrev.124.1866', '10.1088/1478-7814/21/1/321', '10.4401/ag-3741', '10.1038/s41598-019-42892-6', '10.1016/s0264-410x(00)00554-5', '10.1029/94eo00895', None, '10.1073/pnas.76.1.106', '10.1073/pnas.1205553109', '10.1109/mpuls.2019.2937244', '10.1126/science.145.3633.667', '10.1111/j.1574-6968.1992.tb05898.x', None, '10.2427/5688', '10.1016/j.immuni.2010.09.017', '10.1103/physreva.97.023411', '10.1007/s10948-008-0433-x', None, None, '12748315', None, '12375809', None, None, None, None, '28450080', None, None, None, '25207059', '24556987', '16227900', None, '10432482', '26175891', None, '23766957', None, None, '25083827', None, '15458581', '18568940', None, None, '27022144', '10647171', None, None, None, '1462166', '11677681', '20279068', None, None, None, '31015566', '11257410', None, '24713892', '85300', '22753471', None, '14163799', '1384602', '10943392', None, '21029963', None, None, None, None, None, None, '6654177', None, None, None, None, None, None, None, None, '4116029', '3948267', None, None, None, '4498171', None, '3678394', 'title=medicine', None, '4109558', None, None, None, None, None, '4821650', None, None, None, None, None, None, None, None, None, None, '6478851', None, None, '3959394', '382885', '3406819', None, None, None, None, None, '3320742', None, None]","[['acta pharmacologica et toxicologica'], ['the mathematics teacher'], ['new england journal of medicine'], ['nature news'], ['clinical cardiology'], ['[[ieee power '], ['nature '], [' epj web of conferences'], ['archéologie médiévale '], ['neurobiology of learning and memory '], ['technology and culture '], ['monatshefte für mathematik und physik '], ['nature'], ['balkan medical journal'], ['proceedings of the national academy of sciences of the united states of america'], ['spine'], ['performance practice review '], ['neuropsychopharmacology'], ['facts'], ['polymer degradation and stability'], ['beilstein journal of nanotechnology'], ['cambridge university press'], ['radiation research'], ['the journal of clinical investigation'], ['proceedings of the royal society of medicine'], ['neurosurgery '], ['endothelium'], ['physical review'], ['new scientist'], ['journal of experimental medicine'], ['spine'], ['physical review'], ['physical review a'], ['the classical world'], ['seminars in oncology '], ['advances in applied microbiology', 'academic press'], ['nature '], ['physical review'], ['proceedings of the physical society of london'], ['annals of geophysics'], ['scientific reports'], ['vaccine'], ['eos'], ['annals of gastroenterology'], ['proceedings of the national academy of sciences of the united states of america'], ['proceedings of the national academy of sciences'], ['ieee pulse'], ['science '], ['fems microbiology immunology'], ['international microbiology'], ['italian journal of public health'], ['immunity '], ['physical review a'], ['journal of superconductivity and novel magnetism']]",37,5,0,208,0,0,264,0.0647985989492119,0.008756567425569177,0.36427320490367776,0.09982486865148861,0.0,0.1733800350262697,54,"['www.congress.gov', 'energy.gov', 'solarsystem.nasa.gov', 'www.house.gov', 'earthobservatory.nasa.gov', 'www.telecomitalia.com', 'www.britannica.com', 'www.britannica.com', 'www.britannica.com', 'books.google.com', 'www.encyclopedia.com', 'www.britannica.com', 'www.britannica.com', 'www.britannica.com', 'www.britannica.com', 'www.britannica.com', 'www.scientificamerican.com', 'www.britannica.com', 'blogs.discovermagazine.com', 'www.britannica.com', 'www.britannica.com', 'www.thepharmaletter.com', 'www.britannica.com', 'www.britannica.com', 'www.britannica.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'www.timeanddate.com', 'books.google.com', 'www.britannica.com', 'www.britannica.com', 'global.britannica.com', 'www.forgottenweapons.com', 'www.britannica.com', 'www.britannica.com', 'books.google.com', 'thatsmaths.com', 'books.google.com', 'www.conserve-energy-future.com', 'www.biography.com', 'www.britannica.com', 'www.britannica.com', 'www.britannica.com', 'www.choraldirectormag.com', 'vocabulary.com', 'books.google.com', 'www.etymonline.com', 'entertainment.howstuffworks.com', 'www.britannica.com', 'st.ilsole24ore.com', 'www.britannica.com', 'www.britannica.com', 'www.britannica.com', 'www.britannica.com', 'www.britannica.com', 'haloneuroblog.wordpress.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'history.com', 'www.britannica.com', 'www.historyofjeans.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'www.britannica.com', 'www.britannica.com', 'ilglobo.com', 'www.britannica.com', 'www.engineair.com', 'www.britannica.com', 'www.ge.com', 'books.google.com', 'books.google.com', 'courses.lumenlearning.com', 'www.bbgusa.com', 'www.britannica.com', 'www.encyclopedia.com', 'www.britannica.com', 'www.britannica.com', 'www.britannica.com', 'www.autonews.com', 'www.inexhibit.com', 'st.ilsole24ore.com', 'books.google.com', 'www.historyhit.com', 'www.britannica.com', 'www.sms-tsunami-warning.com', 'universityequipe.com', 'www.oldcalculatormuseum.com', 'www.encyclopedia.com', 'www.ilsole24ore.com', 'www.gene.com', 'www.britannica.com', 'www.britannica.com', 'www.britannica.com', 'www.the-scientist.com', 'britannica.com', 'www.classicfm.com', 'www.britannica.com', 'www.britannica.com', 'www.britannica.com', 'faxauthority.com', 'books.google.com', 'materbi.com', 'www.britannica.com', 'www.smithsonianmag.com', 'www.airwaysmuseum.com', 'www.britannica.com', 'www.forbes.com', 'www.britannica.com', 'www.britannica.com', 'www.etymonline.com', 'www.britannica.com', 'bioplasticsnews.com', 'www.britannica.com', 'www.britannica.com', 'www.britannica.com', 'www.britannica.com', 'www.britannica.com', 'linguaggio-macchina.blogspot.com', 'www.castingarea.com', 'www.britannica.com', 'global.britannica.com', 'www.curtamania.com', 'www.oldcalculatormuseum.com', 'newscientist.com', 'www.intel4004.com', 'www.nytimes.com', 'www.britannica.com', 'www.worldatlas.com', 'historyten.com', 'www.britannica.com', 'd-shape.com', 'www.castlesandmanorhouses.com', 'encyclopedia.com', 'about.com', 'www.britannica.com', 'www.museonicolis.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'revivaler.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'encyclopedia.com', 'blog.cheaperthandirt.com', 'www.britannica.com', 'www.engineair.com', 'www.britannica.com', 'www.etymonline.com', 'worldwide.espacenet.com', 'www.britannica.com', 'books.google.com', 'targetitalianideas.com', 'www.britannica.com', 'www.britannica.com', 'www.britannica.com', 'www.britannica.com', 'www.britannica.com', 'www.britannica.com', 'www.britannica.com', 'www.britannica.com', 'www.britannica.com', 'money4u.tripod.com', 'www.britannica.com', 'www.italymagazine.com', 'www.etymonline.com', 'courses.lumenlearning.com', 'patents.justia.com', 'www.britannica.com', 'books.google.com', 'www.smithsonianmag.com', 'europeanconservative.com', 'encyclopedia.com', 'books.google.com', 'www.whonamedit.com', 'www.britannica.com', 'books.google.com', 'www.smithsonianmag.com', 'europeanconservative.com', 'www.telecomitalia.com', 'www.britannica.com', 'intel4004.com', 'www.sciencedaily.com', 'www.britannica.com', 'www.worldatlas.com', 'www.britannica.com', 'onlineeducation.com', 'www.thecollector.com', 'www.britannica.com', 'www.britannica.com', 'www.barcelonayellow.com', 'books.google.com', 'www.topuniversities.com', 'violacentral.com', 'www.britannica.com', 'www.britannica.com', 'www.britannica.com', 'augustobissiri.wordpress.com', 'www.enel.com', 'www.britannica.com', 'books.google.com', 'www.mentalfloss.com', 'newatlas.com', 'www.com', 'nobelprize.org', 'saemobilus.sae.org', 'humanprogress.org', 'www.sciencemag.org', 'collections.nmmusd.org', 'www.famousscientists.org', 'www.iop.org', 'www.edge.org', 'www.nmspacemuseum.org', 'www.internationalpasta.org', 'nobelprize.org', 'www.aacr.org', 'www.orpheon.org', 'www.pbs.org', 'had.aas.org', 'www.msichicago.org', 'www.rasch.org', 'fas.org', 'www.positiveatheism.org', 'www.museoscienza.org', 'edisontechcenter.org', 'nfcnearfieldcommunication.org', 'www.wqxr.org', 'en.irefeurope.org', 'historylists.org', 'rbi.org', 'www.sciencemag.org', 'www.w3.org', 'nobelprize.org', 'www.wqxr.org', 'archive.rubicon-foundation.org', 'museocasertaolivetti.altervista.org', 'edge.org', 'periodic-table.org', 'phys.org', 'museocasertaolivetti.altervista.org', 'phys.org', ['acta pharmacologica et toxicologica'], ['the mathematics teacher'], ['new england journal of medicine'], ['nature news'], ['clinical cardiology'], ['[[ieee power '], ['nature '], [' epj web of conferences'], ['archéologie médiévale '], ['neurobiology of learning and memory '], ['technology and culture '], ['monatshefte für mathematik und physik '], ['nature'], ['balkan medical journal'], ['proceedings of the national academy of sciences of the united states of america'], ['spine'], ['performance practice review '], ['neuropsychopharmacology'], ['facts'], ['polymer degradation and stability'], ['beilstein journal of nanotechnology'], ['cambridge university press'], ['radiation research'], ['the journal of clinical investigation'], ['proceedings of the royal society of medicine'], ['neurosurgery '], ['endothelium'], ['physical review'], ['new scientist'], ['journal of experimental medicine'], ['spine'], ['physical review'], ['physical review a'], ['the classical world'], ['seminars in oncology '], ['advances in applied microbiology', 'academic press'], ['nature '], ['physical review'], ['proceedings of the physical society of london'], ['annals of geophysics'], ['scientific reports'], ['vaccine'], ['eos'], ['annals of gastroenterology'], ['proceedings of the national academy of sciences of the united states of america'], ['proceedings of the national academy of sciences'], ['ieee pulse'], ['science '], ['fems microbiology immunology'], ['international microbiology'], ['italian journal of public health'], ['immunity '], ['physical review a'], ['journal of superconductivity and novel magnetism']]",25829048,Allow all users (no expiry set),240607,16 January 2010,Colonel Warden ,1575,1,2010-01-16,2010-01,2010
507,507,Stonehaven,https://en.wikipedia.org/wiki/Stonehaven,52,0,[],[],4,5,0,6,0,0,37,0.07692307692307693,0.09615384615384616,0.11538461538461539,0.0,0.0,0.17307692307692307,0,"['www.aberdeenshire.gov', 'www.scotlandscensus.gov', 'www.aberdeenshire.gov', 'www.aberdeenshire.gov', 'www.aberdeenshire.gov', 'www.google.com', 'www.fishandchipawards.com', 'www.stunningstonehaven.com', 'www.bbc.com', 'www.heraldscotland.com', 'historic-uk.com', 'journals.socantscot.org', 'www.robertburns.org', 'www.parkrun.org', 'www.warmemorialsonline.org']",156609,Allow all users (no expiry set),33250,10 December 2002,Taras ,653,0,2002-12-10,2002-12,2002
508,508,Rimini,https://en.wikipedia.org/wiki/Rimini,69,1,[],[],0,0,0,17,0,0,51,0.0,0.0,0.2463768115942029,0.014492753623188406,0.0,0.014492753623188406,0,"['www.com', 'www.world-guides.com', 'www.installation-international.com', 'www.com', 'www.com', 'www.ilponte.com', 'statistica.com', 'www.world-guides.com', 'statistica.com', 'www.com', 'www.com', 'www.com', 'www.com', 'www.com', 'it.scribd.com', 'www.britannica.com', 'www.com']",80351,Allow all users (no expiry set),77538,4 September 2002,80.3.160.5 ,984,1,2002-09-04,2002-09,2002
509,509,Aqaba,https://en.wikipedia.org/wiki/Aqaba,82,1,"['10.1023/a:1021196800473', None, None]",[['geojournal']],6,7,0,36,0,0,32,0.07317073170731707,0.08536585365853659,0.43902439024390244,0.012195121951219513,0.0,0.17073170731707318,1,"['www.kinghussein.gov', 'kinghussein.gov', 'nabeul.gov', 'www.dos.gov', 'www.dos.gov', 'www.gov', 'www.nerc.gov', 'books.google.com', 'gcmap.com', 'www.jordantimes.com', 'www.oxfordbusinessgroup.com', 'www.alghad.com', 'www.jpost.com', 'www.addustour.com', 'www.jordantimes.com', 'www.jordantimes.com', 'www.alrai.com', 'books.google.com', 'books.google.com', 'arabiansupplychain.com', 'ynetnews.com', 'books.google.com', 'books.google.com', 'www.yourmiddleeast.com', 'books.google.com', 'jordantimes.com', 'haaretz.com', 'reuters.com', 'addustour.com', 'aqabazone.com', 'www.guinnessworldrecords.com', 'www.addustour.com', 'ynetnews.com', 'www.theworldfolio.com', 'books.google.com', 'www.zawya.com', 'books.google.com', 'www.alghad.com', 'aqabazone.com', 'storymaps.arcgis.com', 'books.google.com', 'www.aqabazone.com', 'www.aqabazone.com', 'lpj.org', 'www.cliohistory.org', 'publications.acorjordan.org', 'www.jreds.org', 'besacenter.org', 'www.jstor.org', ['geojournal']]",328399,Allow all users (no expiry set),69997,27 September 2003,Menchi ,1141,2,2003-09-27,2003-09,2003
510,510,Culture of Rome,https://en.wikipedia.org/wiki/Culture_of_Rome,24,1,"['10.1017/s0009840x00221331', None, None]",[['the classical review ']],3,0,0,7,0,0,13,0.125,0.0,0.2916666666666667,0.041666666666666664,0.0,0.16666666666666666,1,"['romefile.com', 'languagemonitor.com', 'about.com', 'languagemonitor.com', 'books.google.com', 'maspostatevilaregina.com', 'auditorium.com', 'romanculture.org', 'www.archaeology.org', 'www.catholic-hierarchy.org', ['the classical review ']]",25917536,Allow all users (no expiry set),37834,23 January 2010,Theologiae ,185,1,2010-01-23,2010-01,2010
511,511,Bruneian Malay people,https://en.wikipedia.org/wiki/Bruneian_Malay_people,12,0,[],[],0,1,0,7,0,0,4,0.0,0.08333333333333333,0.5833333333333334,0.0,0.0,0.08333333333333333,0,"['www.sabah.gov', 'www.bt.com', 'books.google.com', 'www.bt.com', 'books.google.com', 'books.google.com', 'www.sinarharian.com', 'books.google.com']",23978002,Allow all users (no expiry set),10772,14 August 2009,XPLUSX619 ,265,0,2009-08-14,2009-08,2009
512,512,Da Nang,https://en.wikipedia.org/wiki/Da_Nang,75,0,[],[],1,18,0,17,0,0,39,0.013333333333333334,0.24,0.22666666666666666,0.0,0.0,0.25333333333333335,0,"['www.gso.gov', 'www.gso.gov', '2009-2017.state.gov', 'www.danang.gov', 'danang.gov', 'www.gso.gov', 'vietnamtourism.gov', 'gso.gov', 'www.danang.gov', 'webarchive.loc.gov', 'www.gso.gov', 'www.danang.gov', 'danang.gov', 'danang.gov', 'www.danang.gov', 'www.gso.gov', 'www.danang.gov', 'danang.gov', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'www.angelfire.com', 'www.vietnam-guide.com', 'vietnamnews.vnagency.com', 'worldportsource.com', 'books.google.com', 'www.ttgasia.com', 'www.the-afc.com', 'www.cnn.com', 'www.the-afc.com', 'www.cruisebe.com', 'www.revistapensamientolibre.com', 'books.google.com', 'books.google.com', 'www.vietnam.campusfrance.org']",425140,Allow all users (no expiry set),73133,22 December 2003,Scythian99 ,1426,4,2003-12-22,2003-12,2003
513,513,Bibliography of encyclopedias,https://en.wikipedia.org/wiki/Bibliography_of_encyclopedias,526,2,"['10.4135/9781412965811', '10.1002/9781444338232', None, None, None, None]","[['[[sage publications'], ['wiley-blackwell']]",11,2,0,98,0,0,413,0.02091254752851711,0.0038022813688212928,0.18631178707224336,0.0038022813688212928,0.0,0.028517110266159697,2,"['www.cwb.gov', 'catalogue.nla.gov', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.oxfordreference.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'play.google.com', 'books.google.com', 'books.google.com', 'play.google.com', 'books.google.com', 'books.google.com', 'www.routledge.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.oxfordreference.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.firstworldwar.com', 'www.splashmaritime.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'flagshipmaritimetraining.com', 'books.google.com', 'bivouac.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'amer.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'hypertextbook.com', 'books.google.com', 'books.google.com', 'pwencycl.kgbudge.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.routledge.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'boatcourse.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'play.google.com', 'books.google.com', 'books.google.com', 'play.google.com', 'maritime.org', 's.org', 'pl.wikisource.org', 'oeis.org', 'www.cambridge.org', 's.org', 'www.gutenberg.czyz.org', 'glossary.ametsoc.org', 'www.faqs.org', 'www.guidetoreference.org', 'www.usni.org', ['[[sage publications'], ['wiley-blackwell']]",37062801,Allow all users (no expiry set),297347,19 September 2012,Dr. Blofeld ,2388,2,2012-09-19,2012-09,2012
514,514,Culture of Odisha,https://en.wikipedia.org/wiki/Culture_of_Odisha,6,0,[],[],0,2,0,3,0,0,1,0.0,0.3333333333333333,0.5,0.0,0.0,0.3333333333333333,0,"['www.orissa.gov', 'www.censusindia.gov', 'odishacinema.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com']",17940124,Require administrator access (no expiry set),26341,14 June 2008,Shyamsunder ,339,0,2008-06-14,2008-06,2008
515,515,Catania,https://en.wikipedia.org/wiki/Catania,94,0,[],[],3,2,0,18,0,0,72,0.031914893617021274,0.02127659574468085,0.19148936170212766,0.0,0.0,0.05319148936170213,0,"['www.hko.gov', 'www.catalog.slsa.sa.gov', 'mythindex.com', 'translate.google.com', 'moovitapp.com', 'www.accademiadicatania.com', 'www.cataniaperte.com', 'moovitapp.com', 'bombesullitalia.blogspot.com', 'tripadvisor.mediaroom.com', 'anpi-lissone.over-blog.com', 'www.com', 'etnavalley.com', 'webcache.googleusercontent.com', 'www.collinsdictionary.com', 'weatherbase.com', 'www.agricolturafinanziamenti.com', 'sacramentoritrovato.com', 'tifosobilanciato.wordpress.com', 'en.oxforddictionaries.com', 'creativecommons.org', 'freaknet.org', 'www.cwgc.org']",44776,Allow all users (no expiry set),79050,18 March 2002,62.98.20.244 ,1861,3,2002-03-18,2002-03,2002
516,516,Elizabeth David,https://en.wikipedia.org/wiki/Elizabeth_David,337,1,[],[],30,0,0,15,0,12,279,0.08902077151335312,0.0,0.04451038575667656,0.002967359050445104,0.0,0.09198813056379822,0,"['www.nytimes.com', 'www.nytimes.com', 'www.oxforddnb.com', 'books.google.com', 'www.penguin.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'shop.royalmail.com', 'www.ukwhoswho.com', 'www.nytimes.com', 'www.nytimes.com', 'books.google.com', 'www.penguin.com', 'www.worldcat.org', 'www.worldcat.org', 'www.worldcat.org', 'blog.english-heritage.org', 'www.worldcat.org', 'www.worldcat.org', 'www.worldcat.org', 'www.worldcat.org', 'www.worldcat.org', 'www.worldcat.org', 'www.worldcat.org', 'www.iwm.org', 'www.worldcat.org', 'www.worldcat.org', 'www.worldcat.org', 'www.worldcat.org', 'www.worldcat.org', 'www.worldcat.org', 'www.worldcat.org', 'www.worldcat.org', 'www.worldcat.org', 'www.worldcat.org', 'www.worldcat.org', 'www.worldcat.org', 'www.worldcat.org', 'www.worldcat.org', 'www.worldcat.org', 'www.worldcat.org', 'www.worldcat.org', 'www.english-heritage.org']",1216438,Allow all users (no expiry set),120947,27 November 2004,Bnathyuw ,676,1,2004-11-27,2004-11,2004
517,517,Culture of Russia,https://en.wikipedia.org/wiki/Culture_of_Russia,239,25,"['10.2307/2493225', '10.1038/ejhg.2017.117', '10.1038/s41566-019-0525-0', '10.2307/3020237', '10.2307/125154', '10.1175/1520-0469(1971)028<0263:slovot>2.0.co;2', '10.1080/00085006.2003.11092333', '10.2307/987741', '10.1098/rsbm.1977.0004', '10.2307/2320506', '10.3366/e096813610800037x', '10.1038/nphoton.2007.34', '10.2307/3000442', '10.2307/990455', '10.2307/25587683', '10.2307/27757115', '10.2307/2708192', '10.2307/125254', '10.2307/125968', '10.1016/j.mayocp.2011.11.003', '10.2307/2491790', '10.1080/00085006.1980.11091635', '10.21273/hortsci.50.6.772', '10.2307/127159', None, '28905876', None, None, None, None, None, None, '11615738', None, None, None, None, None, None, None, None, None, None, '22212977', None, None, None, None, None, '5602018', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, '3498096', None, None, None, None]","[['[[slavic review'], ['[[european journal of human genetics'], ['[[nature photonics'], ['[[the slavonic and east european review', '[[cambridge university press'], ['[[wiley ', '[[the russian review'], ['[[academy of sciences of the soviet union', 'journal of the atmospheric sciences'], ['[[canadian slavonic papers'], ['[[journal of the society of architectural historians'], ['[[biographical memoirs of fellows of the royal society'], ['[[taylor ', '[[the american mathematical monthly'], ['[[translation and literature', '[[edinburgh university press'], ['[[nature photonics'], ['[[slavic review', '[[cambridge university press'], ['[[university of california press', '[[journal of the society of architectural historians'], ['the art world'], ['[[university of california press', '[[chymia'], ['[[university of pennsylvania press', '[[journal of the history of ideas'], ['[[the russian review', '[[wiley '], ['[[the russian review', '[[wiley '], ['mayo clinic proceedings '], ['the american slavic and east european review ', '[[association for slavic'], ['[[canadian slavonic papers'], ['hortscience'], ['[[the russian review']]",17,8,0,81,0,7,101,0.07112970711297072,0.03347280334728033,0.3389121338912134,0.10460251046025104,0.0,0.20920502092050208,24,"['2001-2009.state.gov', 'ach.gov', 'history.nasa.gov', 'solarsystem.nasa.gov', 'history.nasa.gov', 'nssdc.gsfc.nasa.gov', 'www.nasa.gov', 'apps.fas.usda.gov', 'www.statista.com', 'www.historytoday.com', 'www.newyorker.com', 'www.discovermagazine.com', 'www.uefa.com', 'www.scimagojr.com', 'www.nytimes.com', 'www.nytimes.com', 'tass.com', 'www.fifa.com', 'books.google.com', 'www.thoughtco.com', 'www.fifa.com', 'www.usatoday.com', 'www.upi.com', 'www.usatoday.com', 'matadornetwork.com', 'www.nytimes.com', 'www.aa.com', 'books.google.com', 'www.rbth.com', 'www.uefa.com', 'www.uefa.com', 'www.statista.com', 'www.bbc.com', 'www.france24.com', 'www.britannica.com', 'mirznanii.com', 'www.themoscowtimes.com', 'www.nybooks.com', 'www.rbth.com', 'filmlinc.com', 'www.rbth.com', 'blogs.transparent.com', 'www.themoscowtimes.com', 'www.geographia.com', 'www.csmonitor.com', 'tass.com', 'encarta.msn.com', 'medium.com', 'www.vox.com', 'www.nytimes.com', 'www.themoscowtimes.com', 'www.euronews.com', 'www.atlasobscura.com', 'www.themoscowtimes.com', 'encarta.msn.com', 'articleswave.com', 'books.google.com', 'www.michigandaily.com', 'slate.com', 'www.britannica.com', 'edition.cnn.com', 'www.history.com', 'www.statista.com', 'www.statista.com', 'www.britannica.com', 'petersburgcity.com', 'www.nytimes.com', 'www.inverse.com', 'qz.com', 'petercioth.medium.com', 'olympics.com', 'www.russia-ic.com', 'nicholaskotar.com', 'www.rbth.com', 'www.rbth.com', 'www.theage.com', 'olympics.com', 'russia-ic.com', 'www.scaruffi.com', 'www.dw.com', 'www.sbs.com', 'www.iihf.com', 'www.dw.com', 'www.rbth.com', 'www.themoscowtimes.com', 'www.forbes.com', 'www.iihf.com', 'www.rlcentre.com', 'www.theatlantic.com', 'medialandscapes.org', 'www.rferl.org', 'www.rferl.org', 'www.russianembassy.org', 'www.npr.org', 'www.jstor.org', 'whc.unesco.org', 'www.npr.org', 'www.rferl.org', 'www.paralympic.org', 'www.rusemb.org', 'www.rferl.org', 'spectrum.ieee.org', 'knightfoundation.org', 'www.bfi.org', 'www.weforum.org', 'gorenka.org', ['[[slavic review'], ['[[european journal of human genetics'], ['[[nature photonics'], ['[[the slavonic and east european review', '[[cambridge university press'], ['[[wiley ', '[[the russian review'], ['[[academy of sciences of the soviet union', 'journal of the atmospheric sciences'], ['[[canadian slavonic papers'], ['[[journal of the society of architectural historians'], ['[[biographical memoirs of fellows of the royal society'], ['[[taylor ', '[[the american mathematical monthly'], ['[[translation and literature', '[[edinburgh university press'], ['[[nature photonics'], ['[[slavic review', '[[cambridge university press'], ['[[university of california press', '[[journal of the society of architectural historians'], ['the art world'], ['[[university of california press', '[[chymia'], ['[[university of pennsylvania press', '[[journal of the history of ideas'], ['[[the russian review', '[[wiley '], ['[[the russian review', '[[wiley '], ['mayo clinic proceedings '], ['the american slavic and east european review ', '[[association for slavic'], ['[[canadian slavonic papers'], ['hortscience'], ['[[the russian review']]",2012490,Allow all users (no expiry set),151796,9 June 2005,Falphin ,2126,10,2005-06-09,2005-06,2005
518,518,Bakewell,https://en.wikipedia.org/wiki/Bakewell,40,0,[],[],2,3,0,7,0,1,27,0.05,0.075,0.175,0.0,0.0,0.125,0,"['www.derbyshiredales.gov', 'www.neighbourhood.statistics.gov', 'www.peakdistrict.gov', 'pitchero.com', 'www.brew-school.com', 'www.newstatesman.com', 'www.pitchero.com', 'rutlandarmsbakewell.com', 'books.google.com', 'britishdelights.com', 'www.oldhousemuseum.org', 'www.bakewellshow.org']",331923,Allow all users (no expiry set),24374,30 September 2003,143.167.21.127 ,628,2,2003-09-30,2003-09,2003
519,519,Corsicans,https://en.wikipedia.org/wiki/Corsicans,33,3,"['10.1038/s41598-019-49901-8', '10.1017/s0021932002002894', '10.1080/03014469600004462', '31537848', '12117210', '8807041', '6753063', None, None]","[['scientific reports'], ['journal of biosocial science'], ['annals of human biology']]",1,0,0,5,0,0,24,0.030303030303030304,0.0,0.15151515151515152,0.09090909090909091,0.0,0.12121212121212122,3,"['maxia-mail.doomby.com', 'books.google.com', 'www.ethnologue.com', 'www.ethnologue.com', 'www.journaldesfemmes.com', 'www.faqs.org', ['scientific reports'], ['journal of biosocial science'], ['annals of human biology']]",3073438,Allow all users (no expiry set),26156,3 November 2005,80.58.192.228 ,522,3,2005-11-03,2005-11,2005
520,520,Palatinate (region),https://en.wikipedia.org/wiki/Palatinate_(region),8,0,[],[],1,0,0,3,0,0,4,0.125,0.0,0.375,0.0,0.0,0.125,0,"['www.britannica.com', 'books.google.com', 'books.google.com', 'www.catholic.org']",38849,Allow all users (no expiry set),23878,11 February 2002,David Parker ,373,0,2002-02-11,2002-02,2002
521,521,Culture of Serbia,https://en.wikipedia.org/wiki/Culture_of_Serbia,55,1,"['0353-5738/2005/0353-57380526065n.pdf', None, None]",[['filozofija i društvo ']],3,0,0,35,0,0,16,0.05454545454545454,0.0,0.6363636363636364,0.01818181818181818,0.0,0.07272727272727272,1,"['books.google.com', 'www.lonelyplanet.com', 'balkaninstitut.com', 'www.rakiabar.com', 'books.google.com', 'books.google.com', 'www.suvenirisrbije.com', 'www.juznevesti.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.festival-cannes.com', 'books.google.com', 'books.google.com', 'espn.com', 'balkaninsight.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'timeshighereducation.com', 'www.crwflags.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.khazars.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'snp.org', 'medialandscapes.org', 'rferl.org', ['filozofija i društvo ']]",2298125,Allow all users (no expiry set),56433,24 July 2005,68.77.145.254 ,696,2,2005-07-24,2005-07,2005
522,522,Sifnos,https://en.wikipedia.org/wiki/Sifnos,24,0,[],[],2,0,0,1,0,0,21,0.08333333333333333,0.0,0.041666666666666664,0.0,0.0,0.08333333333333333,0,"['books.google.com', 'www.stoa.org', 'www.therafoundation.org']",1539931,Allow all users (no expiry set),14358,24 February 2005,62.38.148.30 ,285,1,2005-02-24,2005-02,2005
523,523,Culture of the United Kingdom,https://en.wikipedia.org/wiki/Culture_of_the_United_Kingdom,387,2,"['10.1080/02614367.2010.541481', '10.1159/000144681', None, '970109', None, None]","[[' leisure studies '], ['acta anatomica']]",23,9,0,69,0,13,271,0.059431524547803614,0.023255813953488372,0.17829457364341086,0.00516795865633075,0.0,0.08785529715762273,2,"['www.dft.gov', 'www.legislation.gov', 'www.direct.gov', 'www.statistics.gov', 'www.ons.gov', 'direct.gov', 'www.legislation.gov', 'www.number10.gov', 'www.legislation.gov', 'books.google.com', 'books.google.com', 'www.knebworthhouse.com', 'www.forbes.com', 'names.com', 'www.huffingtonpost.com', 'prideofbritain.com', 'rankings.ft.com', 'www.slate.com', 'copyrighthistory.com', 'www.usatoday.com', 'www.grin.com', 'www.historicfood.com', 'uk.reuters.com', 'www.sesponsorshipgroup.com', 'www.theage.com', 'www.oldmagazinearticles.com', 'books.google.com', 'www.bbc.com', 'www.ft.com', 'books.google.com', 'www.theaustralian.com', 'www.ruleshistory.com', 'www.publishersweekly.com', 'www.ipsos-mori.com', 'homecooking.about.com', 'emotionscards.com', 'books.google.com', 'www.britannica.com', 'edition.cnn.com', 'www.pgatour.com', 'www.nytimes.com', 'www.huffingtonpost.com', 'www.washingtonpost.com', 'www.rolls-roycemotorcars.com', 'www.statista.com', 'fifa.com', 'britannica.com', 'spyhunter007.com', 'tussauds.com', 'www.tennisfame.com', 'www.itv.com', 'www.awardsdaily.com', 'www.heritagebritain.com', 'slate.com', 'www.newsweek.com', 'uefa.com', 'theconversation.com', 'www.britishfashioncouncil.com', 'www.thelondonnottinghillcarnival.com', 'www.itftennis.com', 'www.britannica.com', 'www.britannica.com', 'www.historyextra.com', 'www.rollingstone.com', 'www.time.com', 'www.farminguk.com', 'www.theage.com', 'www.statista.com', 'www.guinnessworldrecords.com', 'postalheritage.wordpress.com', 'www.nytimes.com', 'magazines.com', 'uk.reuters.com', 'books.google.com', 'edition.cnn.com', 'edition.cnn.com', 'www.economist.com', 'www.rampantscotland.com', 'www.english-heritage.org', 'www.ukflavourassociation.org', 'www.gutenberg.org', 'www.the-kennel-club.org', 'olympic.org', 'www.thekennelclub.org', 'britishmuseum.org', 'npg.org', 'www.oldroyalnavalcollege.org', 'dogpages.org', 'www.flaginstitute.org', 'phrases.org', 'www.ymca.org', 'sequart.org', 'scouts.org', 'abbey.org', 'www.scottishtartans.org', 'www.brc.org', 'www.llgc.org', 'www.westminster-abbey.org', 'www.greetingcardassociation.org', 'portal.unesco.org', 'www.jstor.org', [' leisure studies '], ['acta anatomica']]",275009,Allow all users (no expiry set),295023,22 July 2003,Lexor ,4442,1,2003-07-22,2003-07,2003
524,524,Aragon,https://en.wikipedia.org/wiki/Aragon,38,0,[],[],2,0,0,9,0,0,27,0.05263157894736842,0.0,0.23684210526315788,0.0,0.0,0.05263157894736842,0,"['www.rsssf.com', 'www.elperiodicodearagon.com', 'books.google.com', 'www.carnavaldebielsa.com', 'eljusticiadearagon.com', 'datosmacro.com', 'edition.cnn.com', 'www.zaragoza-pirineos2022.com', 'www.elperiodicodearagon.com', 'hdi.globaldatalab.org', 'guara.org']",39443,Allow all users (no expiry set),87755,25 February 2002,David Parker ,1727,2,2002-02-25,2002-02,2002
525,525,Djibouti (city),https://en.wikipedia.org/wiki/Djibouti_(city),40,1,"['10.1080/09397140.2007.10638246', None, None]",[['zoology in the middle east']],5,5,0,9,0,0,20,0.125,0.125,0.225,0.025,0.0,0.275,1,"['www.diyanet.gov', 'addisababa.gov', 'www.weather.gov', 'ftp.atdd.noaa.gov', 'www.cia.gov', 'www.ethnologue.com', 'www.djiboutiairlines.com', 'www.ft.com', 'www.weather-atlas.com', 'djiboutinvest.com', 'www.britannica.com', 'www.washingtonpost.com', 'www.businessinsider.com', 'www.twincities.com', 'hdi.globaldatalab.org', 'www.aaeafrica.org', 'www.comesaria.org', 'www.jstor.org', 'catholic-hierarchy.org', ['zoology in the middle east']]",920729,Allow all users (no expiry set),56191,22 August 2004,WisDom-UK ,1626,0,2004-08-22,2004-08,2004
526,526,Lorraine,https://en.wikipedia.org/wiki/Lorraine,13,0,[],[],0,1,0,1,0,0,11,0.0,0.07692307692307693,0.07692307692307693,0.0,0.0,0.07692307692307693,0,"['minerals.usgs.gov', 'www.lorraineaucoeur.com']",2393620,Allow all users (no expiry set),29749,6 August 2005,Hardouin ,829,0,2005-08-06,2005-08,2005
527,527,Metz,https://en.wikipedia.org/wiki/Metz,186,0,[],[],5,0,0,36,0,0,145,0.026881720430107527,0.0,0.1935483870967742,0.0,0.0,0.026881720430107527,0,"['www.youtube.com', 'www.moselle-tourisme.com', 'www.architecture.com', 'www.youtube.com', 'www.completefrance.com', 'www.fcmetz.com', 'www.meteofrance.com', 'marcmetzmoselle.eklablog.com', 'www.youtube.com', 'www.youtube.com', 'www.lestrinitaires.com', 'meteofrance.com', 'www.tribu.com', 'www.metz-handball.com', 'www.noel-a-metz.com', 'www.shanghairanking.com', 'www.youtube.com', 'www.atpworldtour.com', 'tcrm-blida.com', 'siteindex.francetoday.com', 'www.pnr-lorraine.com', 'www.citadelle-metz.com', 'www.metz-handball.com', 'www.youtube.com', 'www.youtube.com', 'meteofrance.com', 'www.moselle-open.com', 'www.dailymotion.com', 'www.youtube.com', 'www.fcmetz.com', 'tout-metz.com', 'www.ilovemetz.com', 'the95thmovie.com', 'weatherspark.com', 'www.youtube.com', 'www.youtube.com', 'www.fraclorraine.org', 'whc.unesco.org', 'www.quattropole.org', 'whc.unesco.org', 'festival-passages.org']",57906,Allow all users (no expiry set),101078,18 June 2002,Sjc ,1852,2,2002-06-18,2002-06,2002
528,528,List of Spanish inventions and discoveries,https://en.wikipedia.org/wiki/List_of_Spanish_inventions_and_discoveries,41,3,"['10.1021/ed052p325.1', '10.1098/rspl.1854.0094', '10.1002/anie.200330074', None, '30163547', '15376297', None, '5180321', None]","[[' journal of chemical education '], ['proceedings of the royal society of london'], [' angewandte chemie international edition']]",4,1,0,10,0,0,23,0.0975609756097561,0.024390243902439025,0.24390243902439024,0.07317073170731707,0.0,0.1951219512195122,3,"['www.nlm.nih.gov', 'ic.galegroup.com', 'www.livescience.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.typicallyspanish.com', 'www.britannica.com', 'www.lowtechmagazine.com', 'global.oup.com', 'books.google.com', 'www.nobelprize.org', 'ieeeghn.org', 'purl.org', 'www.sfn.org', [' journal of chemical education '], ['proceedings of the royal society of london'], [' angewandte chemie international edition']]",42504960,Allow all users (no expiry set),34852,16 April 2014,Ciudadano001 ,275,0,2014-04-16,2014-04,2014
529,529,Galician culture,https://en.wikipedia.org/wiki/Galician_culture,3,0,[],[],0,0,0,2,0,0,1,0.0,0.0,0.6666666666666666,0.0,0.0,0.0,0,"['maketon.com', 'elprogreso.galiciae.com']",36154048,Allow all users (no expiry set),14809,15 June 2012,Alexander Vigo ,51,0,2012-06-15,2012-06,2012
530,530,Khuzestan province,https://en.wikipedia.org/wiki/Khuzestan_province,42,0,[],[],5,1,0,9,0,0,27,0.11904761904761904,0.023809523809523808,0.21428571428571427,0.0,0.0,0.14285714285714285,0,"['www.eia.gov', 'www.janes.com', 'bbcpersian.com', 'kojaro.com', 'www.iranchamber.com', 'books.google.com', 'statoids.com', 'aparat.com', 'parsine.com', 'iranica.com', 'hdi.globaldatalab.org', 'www.amar.org', 'www.iftiz.org', 'www.sci.org', 'amar.org']",448079,Allow all users (no expiry set),52590,30 January 2004,Morwen ,1665,3,2004-01-30,2004-01,2004
531,531,Tourism in the Basque Autonomous Community,https://en.wikipedia.org/wiki/Tourism_in_the_Basque_Autonomous_Community,20,0,[],[],1,0,0,4,0,0,15,0.05,0.0,0.2,0.0,0.0,0.05,0,"['www.tripadvisor.com', 'eitb.com', 'www.surfingeuskadi.com', 'sallybernstein.com', 'vitoria-gasteiz.org']",33516239,Allow all users (no expiry set),22683,24 October 2011,Saboreala ,78,0,2011-10-24,2011-10,2011
532,532,Aleppo,https://en.wikipedia.org/wiki/Aleppo,191,3,"['10.1093/ehr/xcv.ccclxxvi.481', '10.1163/15700658-bja10030', '10.1080/00291463.1972.11675812', None, None, None, None, None, None]","[['[[the english historical review'], ['journal of early modern history '], ['nordisk psykologi']]",22,1,0,95,0,3,67,0.11518324607329843,0.005235602094240838,0.4973821989528796,0.015706806282722512,0.0,0.13612565445026178,3,"['ftp.atdd.noaa.gov', 'almaany.com', 'books.google.com', 'books.google.com', 'www.trtworld.com', 'www.reuters.com', 'www.cbsnews.com', 'worldpopulationreview.com', 'armenianweekly.com', 'madinatuna.com', 'www.britannica.com', 'www.worldstadiums.com', 'www.nytimes.com', 'www.cpamedia.com', 'books.google.com', 'syrcata.com', 'books.google.com', 'everything2.com', 'www.almasdarnews.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.nytimes.com', 'emirates247.com', 'books.google.com', 'kyivpost.com', 'imageusa.com', 'www.heraldsun.com', 'aksalser.com', 'books.google.com', 'brill.com', 'books.google.com', 'www.isalep.com', 'dp-news.com', 'heartoforient.blogspot.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'madinatuna.com', 'www.almasdarnews.com', 'www.reuters.com', 'www.nytimes.com', 'brill.com', 'books.google.com', 'www.reuters.com', 'syria-news.com', 'middleeast.com', 'www.imsoblesseddaily.com', 'edition.cnn.com', 'apnews.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.ursoap.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'aliqtisadi.com', 'www.reuters.com', 'www.dailystar.com', 'syrianhistory.com', 'books.google.com', 'books.google.com', 'brill.com', 'www.ibtimes.com', 'www.irishtimes.com', 'books.google.com', 'www.dp-news.com', 'books.google.com', 'forward.com', 'www.aljazeera.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.haaretz.com', 'books.google.com', 'books.google.com', 'www.dnnar.com', 'www.bbc.com', 'www.dailysabah.com', 'books.google.com', 'en.oxforddictionaries.com', 'www.syriasteps.com', 'www.newyorker.com', 'www.nytimes.com', 'www.aksalser.com', 'www.syria-news.com', 'www.almasdarnews.com', 'brill.com', 'panoramaline.com', 'edition.cnn.com', 'aina.org', 'www.udp-aleppo.org', 'www.worldheritagesite.org', 'www.terezia.org', 'www.npr.org', 'www.aladeyat.org', 'www.cbssyr.org', 'data.un.org', 'archnet.org', 'whc.unesco.org', 'syriacpatriarchate.org', 'www.syria.strabon.org', 'www.syriatourism.org', 'en.unesco.org', 'www.thirdrva.org', 'www.cbssyr.org', 'carnegie-mec.org', 'whc.unesco.org', 'www.cbssyr.org', 'www.terezia.org', 'www.cbssyr.org', 'www.cambridge.org', ['[[the english historical review'], ['journal of early modern history '], ['nordisk psykologi']]",159244,Allow all users (no expiry set),164808,18 December 2002,62.253.64.7 ,4238,15,2002-12-18,2002-12,2002
533,533,Culture of Brisbane,https://en.wikipedia.org/wiki/Culture_of_Brisbane,12,0,[],[],0,0,0,11,0,0,1,0.0,0.0,0.9166666666666666,0.0,0.0,0.0,0,"['www.zomato.com', 'www.zomato.com', 'www.zomato.com', 'publicartwork.jsadigital.com', 'www.zomato.com', 'www.visitbrisbane.com', 'www.zomato.com', 'www.zomato.com', 'www.zomato.com', 'www.zomato.com', '2015.buddhabirthdayfestival.com']",3748328,Allow all users (no expiry set),19441,17 January 2006,CJ ,303,0,2006-01-17,2006-01,2006
534,534,Haryanvi people,https://en.wikipedia.org/wiki/Haryanvi_people,17,0,[],[],1,1,0,12,0,0,3,0.058823529411764705,0.058823529411764705,0.7058823529411765,0.0,0.0,0.11764705882352941,0,"['csharyana.gov', 'books.google.com', 'www.expressindia.com', 'iitd.ac.com', 'books.google.com', 'www.hindu.com', 'www.livemint.com', 'www.pressreader.com', 'articles.timesofindia.indiatimes.com', 'www.tribuneindia.com', 'books.google.com', 'books.google.com', 'www.tribuneindia.com', 'multitree.org']",63497599,Allow all users (no expiry set),13731,28 March 2020,Dev0745 ,160,2,2020-03-28,2020-03,2020
535,535,History of the Jews in Los Angeles,https://en.wikipedia.org/wiki/History_of_the_Jews_in_Los_Angeles,62,0,[],[],10,0,0,39,0,0,14,0.16129032258064516,0.0,0.6290322580645161,0.0,0.0,0.16129032258064516,0,"['articles.latimes.com', 'lubavitch.com', 'www.washingtonpost.com', 'haruth.com', 'books.google.com', 'www.dailynews.com', 'jewishexponent.com', 'articles.latimes.com', 'articles.latimes.com', 'nl.newsbank.com', 'articles.latimes.com', 'www.latimes.com', 'www.latimes.com', 'www.latimes.com', 'newsok.com', 'business.highbeam.com', 'www.ateretisrael.com', 'books.google.com', 'www.multichannel.com', 'articles.latimes.com', 'www.laweekly.com', 'chabad.com', 'books.google.com', 'www.daytrippertours.com', 'www.latimes.com', 'www.dailynews.com', 'books.google.com', 'www.wmagazine.com', 'articles.latimes.com', 'rogerebert.com', 'www.haaretz.com', 'www.chabaducla.com', 'jewishjournal.com', 'www.jewishjournal.com', 'jewishjournal.com', 'jewishjournal.com', 'articles.latimes.com', 'www.latimes.com', 'articles.latimes.com', 'www.jewishla.org', 'iajf.org', 'newsreel.org', 'www.jewishdatabank.org', 'perspectives.ajsnet.org', 'www.jewishla.org', 'www.shturem.org', 'chabad.org', 'dbs.bh.org', 'www.jewishfilm.org']",42358585,Allow all users (no expiry set),56567,31 March 2014,WhisperToMe ,319,0,2014-03-31,2014-03,2014
536,536,Diyarbakır,https://en.wikipedia.org/wiki/Diyarbak%C4%B1r,98,8,"['10.1093/acref/9780198662778.001.0001', '10.1017/s0896634600004180', '10.1353/anq.2017.0004', '10.1525/jsah.2014.73.4.507', '10.1017/s0010417512000400', '10.1080/00263209608701112', '10.23976/smep.2014008', None, None, None, None, None, None, None, None, None, None, None, None, None, None]","[['oxford university press'], ['new perspectives on turkey'], ['anthropological quarterly'], ['journal of the society of architectural historians'], ['comparative studies in society and history'], ['middle eastern studies'], ['singapore middle east papers']]",17,3,0,33,0,0,37,0.17346938775510204,0.030612244897959183,0.336734693877551,0.08163265306122448,0.0,0.2857142857142857,7,"['www.mgm.gov', 'diyarbakir.meb.gov', 'arastirma.tarimorman.gov', 'www.al-monitor.com', 'ahvalnews.com', 'books.google.com', 'sabah.com', 'westarmgen.weebly.com', 'www.alevinet.com', 'romeartlover.tripod.com', 'www.nytimes.com', 'www.hurriyetdailynews.com', 'www.radikal.com', 'www.milliyet.com', 'books.google.com', 'www.turkishairlines.com', 'www.almasdarnews.com', 'books.google.com', 'yektauzunoglu.com', 'www.aljazeera.com', 'www.haberturk.com', 'www.ensonhaber.com', 'www.suryaniler.com', 'www.lonelyplanet.com', 'secim.haberler.com', 'www.hurriyetdailynews.com', 'www.agos.com', 'referenceworks.brillonline.com', 'www.euronews.com', 'www.hurriyetdailynews.com', 'books.google.com', 'www.diyarbakirsoz.com', 'books.google.com', 'books.google.com', 'www.france24.com', 'www.bbc.com', 'escholarship.org', 'www.wdl.org', 'whc.unesco.org', 'www.arkeologlardernegist.org', 'www.bianet.org', 'www.wdl.org', 'www.worldcat.org', 'www.lalishduhok.org', 'www.wdl.org', 'www.wdl.org', 'www.wdl.org', 'www.worldcat.org', 'worldcat.org', 'www.hrw.org', 'www.worldcat.org', 'www.worldcat.org', 'sedra.bethmardutho.org', ['oxford university press'], ['new perspectives on turkey'], ['anthropological quarterly'], ['journal of the society of architectural historians'], ['comparative studies in society and history'], ['middle eastern studies'], ['singapore middle east papers']]",642286,Allow all users (no expiry set),66273,8 May 2004,81.215.13.201 ,2082,8,2004-05-08,2004-05,2004
537,537,Rastoke,https://en.wikipedia.org/wiki/Rastoke,0,0,[],[],0,0,0,0,0,0,0,,,,,,,0,[],2787544,Allow all users (no expiry set),14960,28 September 2005,Maestral ,123,0,2005-09-28,2005-09,2005
538,538,Northern England,https://en.wikipedia.org/wiki/Northern_England,361,3,"['10.1002/joc.1276', '10.2307/213484', '10.1080/14797585.2015.1134056', None, None, None, None, None, None]","[['international journal of climatology'], ['geographical review'], ['journal for cultural research']]",32,35,0,74,0,22,196,0.0886426592797784,0.09695290858725762,0.20498614958448755,0.008310249307479225,0.0,0.19390581717451524,3,"['webarchive.nationalarchives.gov', 'www.metoffice.gov', 'www.gov', 'www.gov', 'www.gov', 'www.gov', 'www.ons.gov', 'www.ons.gov', 'www.ons.gov', 'www.ons.gov', 'www.gov', 'www.metoffice.gov', 'www.ons.gov', 'www.metoffice.gov', 'www.leeds.gov', 'www.ons.gov', 'www.gov', 'www.ons.gov', 'www.lakedistrict.gov', 'www.ons.gov', 'www.ons.gov', 'www.gov', 'www.ons.gov', 'www.ons.gov', 'webarchive.nationalarchives.gov', 'statistics.gov', 'www.metoffice.gov', 'www.ons.gov', 'www.gov', 'www.gov', 'www.ons.gov', 'www.ons.gov', 'www.gov', 'www.gov', 'www.metoffice.gov', 'www.itv.com', 'www.ft.com', 'www.transportforthenorth.com', 'www.skysports.com', 'www.buzzfeed.com', 'www.historytoday.com', 'books.google.com', 'tech.newstatesman.com', 'www.visitengland.com', 'www.fifa.com', 'www.ft.com', 'www.reuters.com', 'books.google.com', 'books.google.com', 'www.citymetric.com', 'www.bbc.com', 'theconversation.com', 'www.ft.com', 'universityhistories.com', 'origin.misc.pagesuite.com', 'thetab.com', 'www.bbc.com', 'www.ft.com', 'www.railjournal.com', 'time.com', 'www.vanityfair.com', 'www.citymetric.com', 'www.englandsimmigrants.com', 'www.newstatesman.com', 'www.bbc.com', 'books.google.com', 'www.newstatesman.com', 'www.transportforthenorth.com', 'www.bbc.com', 'www.bbc.com', 'www.dazeddigital.com', 'www.focus-economics.com', 'www.newstatesman.com', 'www.citymetric.com', 'www.newstatesman.com', 'books.google.com', 'www.ft.com', 'books.google.com', 'www.jewishencyclopedia.com', 'books.google.com', 'www.citymetric.com', 'www.economist.com', 'www.britishelectionstudy.com', 'books.google.com', 'www.buzzfeed.com', 'www.bbc.com', 'www.bbc.com', 'www.economist.com', 'www.bbc.com', 'carlscam.com', 'www.bbc.com', 'www.radiotimes.com', 'www.bbc.com', 'www.bbc.com', 'www.britishheritage.com', 'www.uktradeinfo.com', 'www.visitengland.com', 'medicalxpress.com', 'www.goldenageofnorthumbria.com', 'www.bbcgoodfood.com', 'www.techradar.com', 'books.google.com', 'www.citymetric.com', 'www.newstatesman.com', 'www.historytoday.com', 'www.citymetric.com', 'books.google.com', 'books.google.com', 'books.google.com', 'bcw-project.org', 'www.liverpoolmuseums.org', 'naturalengland.org', 'mosques.muslimsinbritain.org', 'mosques.muslimsinbritain.org', 'www.n8research.org', 'www.ippr.org', 'www.britishcouncil.org', 'www.cbi.org', 'www.ippr.org', 'www.electoralcommission.org', 'www.webarchive.org', 'www.r-c.org', 'lindisfarne.org', 'www.visitbritain.org', 'waterwise.org', 'research.historicengland.org', 'www.yorkshiredialectsociety.org', 'bcw-project.org', 'www.northumbriana.org', 'www.fao.org', 'www.greatrun.org', 'www.ehs.org', 'www.visitbritain.org', 'humanism.org', 'www.dockmuseum.org', 'canalrivertrust.org', 'waterwise.org', 'www.railnorth.org', 'www.newsworks.org', 'search.electoralcommission.org', 'www.ippr.org', ['international journal of climatology'], ['geographical review'], ['journal for cultural research']]",714694,Allow all users (no expiry set),232949,10 June 2004,Morwen ,2318,1,2004-06-10,2004-06,2004
539,539,List of Austrian inventions and discoveries,https://en.wikipedia.org/wiki/List_of_Austrian_inventions_and_discoveries,1,0,[],[],0,0,0,0,0,0,1,0.0,0.0,0.0,0.0,0.0,0.0,0,[],39265475,Allow all users (no expiry set),3581,30 April 2013,WienaBerlina ,58,0,2013-04-30,2013-04,2013
540,540,Syldavia,https://en.wikipedia.org/wiki/Syldavia,9,0,[],[],0,0,0,3,0,0,6,0.0,0.0,0.3333333333333333,0.0,0.0,0.0,0,"['www.google.com', 'www.google.com', 'books.google.com']",54552,Allow all users (no expiry set),19774,1 June 2002,PierreAbbat ,667,0,2002-06-01,2002-06,2002
541,541,Cham Albanians,https://en.wikipedia.org/wiki/Cham_Albanians,295,6,"['10.4000/ejts.4444', '10.1525/ae.1999.26.1.196', '10.12681/eadd/33128', '10.1525/ah.2005.79.3.321', '10.12681/eadd/17487', '10.2307/1785338', None, None, None, None, None, None, None, None, None, None, None, None]","[['european journal of turkish studies. social sciences on contemporary turkey', 'european journal of turkish studies'], ['american ethnologist'], ['[[democritus university of thrace'], ['department of history', 'agricultural history'], ['panteion university of social and political sciences'], ['the geographical journal']]",10,1,0,105,0,0,173,0.03389830508474576,0.003389830508474576,0.3559322033898305,0.020338983050847456,0.0,0.0576271186440678,6,"['www.qpz.gov', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.pdi-al.com', 'books.google.com', 'books.google.com', 'vasiltole.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'adherents.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.pdu-al.com', 'books.google.com', 'katoci.blogspot.com', 'vasiltole.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'chameriaorganization.blogspot.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.ceeol.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thefreedictionary.com', 'books.google.com', 'books.google.com', 'www.ceeol.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.balkaninsight.com', 'www.ceeol.com', 'books.google.com', 'books.google.com', 'www.geocities.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.milliyet.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.ethnologue.com', 'www.ceeol.com', 'books.google.com', 'books.google.com', 'books.google.com', 'krahuishqiponjes.blogspot.com', 'books.google.com', 'adherents.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.ceeol.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.chameriaassociation.org', 'ejts.revues.org', 'www.cec.org', 'www.rferl.org', 'www.imir-bg.org', 'imir-bg.org', 'cameriainstitute.org', 'www.farsarotul.org', 'balkanologie.revues.org', 'www.eens.org', ['european journal of turkish studies. social sciences on contemporary turkey', 'european journal of turkish studies'], ['american ethnologist'], ['[[democritus university of thrace'], ['department of history', 'agricultural history'], ['panteion university of social and political sciences'], ['the geographical journal']]",309105,Allow all users (no expiry set),256721,1 September 2003,Wik ,2983,0,2003-09-01,2003-09,2003
542,542,Culture of Poland,https://en.wikipedia.org/wiki/Culture_of_Poland,11,0,[],[],0,1,0,0,0,0,10,0.0,0.09090909090909091,0.0,0.0,0.0,0.09090909090909091,0,['poland.gov'],1626892,Allow all users (no expiry set),34103,20 March 2005,Piotrus ,836,4,2005-03-20,2005-03,2005
543,543,Adana,https://en.wikipedia.org/wiki/Adana,148,2,"['10.1186/bf03352554', '10.1163/15700658-bja10030', None, None, None, None]","[['earth planets space '], ['journal of early modern history ']]",22,19,0,60,0,0,45,0.14864864864864866,0.12837837837837837,0.40540540540540543,0.013513513513513514,0.0,0.2905405405405405,2,"['www.ogm-adanaobm.gov', 'adana.meb.gov', 'www.tbmm.gov', 'www.adanaozelidare.gov', 'biruni.tuik.gov', 'adana.gov', 'www.ogm-adanaobm.gov', 'www.tbmm.gov', 'www.adanadt.gov', 'www.adanakultur.gov', 'www.adanakutup.gov', 'www.mgm.gov', 'adana.ktb.gov', 'thf.gov', 'adana-bld.gov', 'adana-bld.gov', 'todd.gov', 'www.dhmi.gov', 'thf.gov', 'www.todor66.com', 'www.agos.com', 'www.mekan360.com', 'karar.com', 'www.adonisistanbul.com', 'www.habername.com', 'www.sabah.com', 'books.google.com', 'www.fdimagazine.com', 'www.radikal.com', 'www.sabah.com', 'gazeteolay.com', 'birdeburadandinleyin.blogspot.com', 'www.kenthaber.com', 'www.sondakika.com', 'spor.haberler.com', 'www.universityworldnews.com', 'www.advansa.com', 'www.agos.com', 'www.adanakentkutuphanesi.com', 'haber.gazetevatan.com', 'cezmiyurtsever.com', 'books.google.com', 'www.flyair.com', 'haber01.com', 'haberler.com', 'gezily.com', 'www.medikalplus.com', 'haberler.com', 'haberler.com', 'www.sabah.com', 'www.bolgegundem.com', 'cnnturk.com', 'haberler.com', 'issuu.com', 'www.kenthaber.com', 'www.kentselhaber.com', 'www.marsangida.com', 'www.hurriyet.com', 'www.tumgazeteler.com', 'www.tuyap.com', 'bourjhammoud.com', 'www.zaman.com', 'haberler.com', 'www.radikal.com', 'www.hyeetch.nareg.com', 'www.haberler.com', 'www.haberler.com', 'books.google.com', 'books.google.com', 'www.adanamedya.com', 'nisandaadanada.com', 'www.dunyagazetesi.com', 'books.google.com', 'haberler.com', 'www.aksiyon.com', 'www.radikal.com', 'www.cukobirlik.com', 'haberler.com', 'www.stargazete.com', 'www.azsam.org', 'tff.org', 'www.imo.org', 'www.anadolukatolikkilisesi.org', 'www.hri.org', 'www.adana-to.org', 'www.adaso.org', 'www.adanatb.org', 'www.iranicaonline.org', 'tvf.org', 'www.worldhistory.org', 'www.adanademirspor.org', 'www.cumder.org', 'www.atonet.org', 'www.worldhistory.org', 'www.turkyaybir.org', 'www.sabancivakfi.org', 'hrantdink.org', 'www.cuktob.org', 'hrantdink.org', 'seyahat.buneki.org', 'sabancivakfi.org', ['earth planets space '], ['journal of early modern history ']]",185243,Allow all users (no expiry set),152694,19 February 2003,Susan Mason ,4755,11,2003-02-19,2003-02,2003
544,544,List of English words of Russian origin,https://en.wikipedia.org/wiki/List_of_English_words_of_Russian_origin,12,0,[],[],0,0,0,3,0,0,9,0.0,0.0,0.25,0.0,0.0,0.0,0,"['www.oed.com', 'www.oed.com', 'observer.com']",402136,Allow all users (no expiry set),68386,15 December 2003,Ilya ,1031,1,2003-12-15,2003-12,2003
545,545,Aksaray,https://en.wikipedia.org/wiki/Aksaray,14,0,[],[],1,4,0,4,0,0,5,0.07142857142857142,0.2857142857142857,0.2857142857142857,0.0,0.0,0.35714285714285715,0,"['data.tuik.gov', 'www.harita.gov', 'aksaray.turizm.gov', 'www.mgm.gov', 'books.google.com', 'bizimil.com', 'www.yenisafak.com', 'www.fallingrain.com', 'icvbbulletin.org']",1651292,Allow all users (no expiry set),24504,26 March 2005,Sezaiata ,416,1,2005-03-26,2005-03,2005
546,546,"Brest, France","https://en.wikipedia.org/wiki/Brest,_France",37,0,[],[],4,2,0,10,0,0,21,0.10810810810810811,0.05405405405405406,0.2702702702702703,0.0,0.0,0.16216216216216217,0,"['ftp.atdd.noaa.gov', 'www.plymouth.gov', 'www.etymonline.com', 'www.avidcruiser.com', 'www.completefrance.com', 'www.railwaygazette.com', 'www.meteofrance.com', 'books.google.com', 'brest.letelegramme.com', 'www.britannica.com', 'www.meteofrance.com', 'edition.cnn.com', 'denversistercities.org', 'upload.wikimedia.org', 'www.ofis-bzh.org', 'nizkor.org']",57912,Allow all users (no expiry set),46562,18 June 2002,Jeronimo ,1099,0,2002-06-18,2002-06,2002
547,547,Culture of South Africa,https://en.wikipedia.org/wiki/Culture_of_South_Africa,27,3,"['10.2989/16073614.2011.633360', '10.1080/02560046.2019.1647256', None, None, None, None]","[['southern african linguistics and applied language studies'], ['critical arts']]",5,0,0,8,0,2,9,0.18518518518518517,0.0,0.2962962962962963,0.1111111111111111,0.0,0.2962962962962963,2,"['books.google.com', 'www.youtube.com', 'findarticles.com', 'www.riaa.com', 'findarticles.com', 'www.news24.com', 'www.news24.com', 'www.youtube.com', 'hdr.undp.org', 'www.actionaid.org', 'teachenglishtoday.org', 'www.sodomylaws.org', 'www.scouting.org', ['southern african linguistics and applied language studies'], ['critical arts']]",364917,Allow all users (no expiry set),33225,12 November 2003,Boffin ,1197,0,2003-11-12,2003-11,2003
548,548,"Rampur, Uttar Pradesh","https://en.wikipedia.org/wiki/Rampur,_Uttar_Pradesh",46,0,[],[],1,4,0,27,0,0,14,0.021739130434782608,0.08695652173913043,0.5869565217391305,0.0,0.0,0.10869565217391304,0,"['pib.gov', 'razalibrary.gov', 'razalibrary.gov', 'censusindia.gov', 'www.amarujala.com', 'www.indiantoners.com', 'www.wheelsindia.com', 'www.indiainfoline.com', 'indianexpress.com', 'www.business-standard.com', 'www.source2update.com', 'www.milligazette.com', 'www.sunwayschool.com', 'whitehallpublicschool.com', 'www.flickr.com', 'www.menthaallied.com', 'radicokhaitan.com', 'amritvichar.com', 'www.dmarampur.com', 'www.nainitaltourism.com', 'hoparoundindia.com', 'gmail.com', 'www.indianexpress.com', 'www.nainitaltourism.com', 'www.ustadrashidkhan.com', 'www.livemint.com', 'india9.com', 'www.thehindu.com', 'www.hoparoundindia.com', 'www.indiablooms.com', 'india9.com', 'stjohntanda.org']",517319,Allow all users (no expiry set),46320,10 March 2004,18.234.1.84 ,1133,2,2004-03-10,2004-03,2004
549,549,Arab culture,https://en.wikipedia.org/wiki/Arab_culture,60,6,"['10.1177/001654929605800102', '10.1080/14616700802337800', '10.1177/1748048506062233', '10.1177/0016549299061001004', '10.1177/1940161208317142', None, None, None, None, None, None, None, None, None, None]","[['international communication gazette'], ['journalism studies'], ['international communication gazette'], ['international communication gazette'], ['the international journal of press']]",2,0,0,21,0,0,31,0.03333333333333333,0.0,0.35,0.1,0.0,0.13333333333333333,5,"['www.youtube.com', 'fifa.com', 'arabmediasociety.com', 'fifa.com', 'www.youtube.com', 'books.google.com', 'jordantimes.com', 'al-bab.com', 'thelede.blogs.nytimes.com', 'www.ikhwanweb.com', 'ourpastimes.com', 'www.aljazeera.com', 'bayt.com', 'www.youtube.com', 'muslimwomeninsports.blogspot.com', 'www.arabmediasociety.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.arabmediasociety.com', 'www.youtube.com', 'fas.org', 'cpj.org', ['international communication gazette'], ['journalism studies'], ['international communication gazette'], ['international communication gazette'], ['the international journal of press']]",4087576,Allow all users (no expiry set),67333,16 February 2006,Marudubshinki ,1080,3,2006-02-16,2006-02,2006
550,550,Culture of Croatia,https://en.wikipedia.org/wiki/Culture_of_Croatia,23,0,[],[],3,0,0,1,0,0,19,0.13043478260869565,0.0,0.043478260869565216,0.0,0.0,0.13043478260869565,0,"['artchive.com', 'faostat.fao.org', 'www.rastko.org', 'www.disabilityartsonline.org']",474950,Allow all users (no expiry set),32210,18 February 2004,Joy ,536,1,2004-02-18,2004-02,2004
551,551,Shiga Prefecture,https://en.wikipedia.org/wiki/Shiga_Prefecture,19,0,[],[],0,0,0,1,0,0,18,0.0,0.0,0.05263157894736842,0.0,0.0,0.0,0,['www.oumiushi.com'],179773,Allow all users (no expiry set),33304,6 February 2003,Synthetik ,481,5,2003-02-06,2003-02,2003
552,552,Gurage people,https://en.wikipedia.org/wiki/Gurage_people,19,0,[],[],1,3,0,1,0,0,14,0.05263157894736842,0.15789473684210525,0.05263157894736842,0.0,0.0,0.21052631578947367,0,"['www.csa.gov', 'www.csa.gov', 'www.csa.gov', 'books.google.com', 'www.worldcat.org']",1619668,Allow all users (no expiry set),16973,18 March 2005,Shiferaw ,1094,3,2005-03-18,2005-03,2005
553,553,Tourism in Finland,https://en.wikipedia.org/wiki/Tourism_in_Finland,35,0,[],[],2,0,0,14,0,0,19,0.05714285714285714,0.0,0.4,0.0,0.0,0.05714285714285714,0,"['saunafromfinland.com', 'www.travelpricewatch.com', 'finlandprices.com', 'www.worldairportawards.com', 'touch.lonelyplanet.com', 'ubs.com', 'misstourist.com', 'theculturetrip.com', 'businesstampere.com', 'travelpricewatch.com', 'www.finlandprices.com', 'www.timeshighereducation.com', 'travelmelodies.com', 'www.spottedbylocals.com', 'www.baltic.org', 'search.isepstudyabroad.org']",159637,Allow all users (no expiry set),23525,19 December 2002,212.59.40.55 ,356,0,2002-12-19,2002-12,2002
554,554,Province of Parma,https://en.wikipedia.org/wiki/Province_of_Parma,1,0,[],[],0,0,0,0,0,0,1,0.0,0.0,0.0,0.0,0.0,0.0,0,[],987110,Allow all users (no expiry set),12093,15 September 2004,Stan Shebs ,158,0,2004-09-15,2004-09,2004
555,555,Póvoa de Varzim,https://en.wikipedia.org/wiki/P%C3%B3voa_de_Varzim,192,0,[],[],7,4,0,19,0,0,162,0.036458333333333336,0.020833333333333332,0.09895833333333333,0.0,0.0,0.057291666666666664,0,"['www.autarquicas2021.mai.gov', 'nasa.gov', 'www.diramb.gov', 'digitarq.dgarq.gov', 'maximusproject.com', 'www.povoadevarzim.com', 'www.correiodabeiraserra.com', 'www.slowfoodfoundation.com', 'www.catholic-forum.com', 'www.povoadevarzim.com', 'www.aeroclubedonorte.com', 'www.golfdigest.com', 'www.lifecooler.com', 'hatcheryinternational.com', 'www.sail-world.com', 'maximusproject.com', 'uk.news.yahoo.com', 'www.newgreenfil.com', 'virtualbooks.terra.com', 'www2.elmundolibro.com', 'www.oceanpd.com', 'www.fpnatacao.com', 'www.povoadevarzim.com', 'www.oecd.org', 'www.profissionaisdoscasinos.org', 'www.portugalpride.org', 'eurekalert.org', 'www.turismoreligioso.org', 'www.fatima.org', 'vialivre.org']",316446,Allow all users (no expiry set),153958,12 September 2003,194.65.14.70 ,2075,2,2003-09-12,2003-09,2003
556,556,Boro culture,https://en.wikipedia.org/wiki/Boro_culture,9,1,"['10.1016/j.dit.2013.09.002', None, None]",[['drug invention today ']],0,1,0,0,0,0,7,0.0,0.1111111111111111,0.0,0.1111111111111111,0.0,0.2222222222222222,1,"['www.udalguri.gov', ['drug invention today ']]",7246558,Allow all users (no expiry set),10177,1 October 2006,Chaipau ,295,0,2006-10-01,2006-10,2006
557,557,Cappadocian Greeks,https://en.wikipedia.org/wiki/Cappadocian_Greeks,119,0,[],[],1,0,0,7,0,0,111,0.008403361344537815,0.0,0.058823529411764705,0.0,0.0,0.008403361344537815,0,"['www.gettyimages.com', 'books.google.com', 'www.khamush.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.hurriyetdailynews.com', 'www.kms.org']",36492342,Allow all users (no expiry set),133303,20 July 2012,Zorlusert ,294,2,2012-07-20,2012-07,2012
558,558,Kayseri,https://en.wikipedia.org/wiki/Kayseri,20,0,[],[],5,1,0,7,0,0,7,0.25,0.05,0.35,0.0,0.0,0.3,0,"['www.mgm.gov', 'www.kayser.com', 'myweather2.com', 'www.scribd.com', 'gezily.com', 'books.google.com', 'www.oxfordreference.com', 'books.google.com', 'www.tff.org', 'esiweb.org', 'www.virtualani.org', 'www.jstor.org', 'www.esiweb.org']",242346,Allow all users (no expiry set),32108,8 June 2003,195.87.131.93 ,1130,2,2003-06-08,2003-06,2003
559,559,Baghdadi Jews,https://en.wikipedia.org/wiki/Baghdadi_Jews,73,3,"['10.1017/s0026749x03004104', '10.1353/sho.0.0213', '10.2307/3622197', None, None, None, None, None, None]","[['modern asian studies'], ['shofar'], ['proceedings of the american academy for jewish research']]",14,1,0,45,0,0,10,0.1917808219178082,0.0136986301369863,0.6164383561643836,0.0410958904109589,0.0,0.2465753424657534,3,"['www.ija.archives.gov', 'issuu.com', 'forward.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.penangjewishcemetery.com', 'books.google.com', 'www.dangoor.com', 'books.google.com', 'books.google.com', 'thejc.com', 'www.openthemagazine.com', 'books.google.com', 'www.myjewishlearning.com', 'books.google.com', 'rangandatta.wordpress.com', 'books.google.com', 'books.google.com', 'books.google.com', 'india.blogs.nytimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'singaporejews.com', 'books.google.com', 'tabletmag.com', 'granta.com', 'india.blogs.nytimes.com', 'books.google.com', 'books.google.com', 'jewsofjava.com', 'referenceworks.brillonline.com', 'books.google.com', 'www.haaretz.com', 'books.google.com', 'issuu.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.jstor.org', 'www.jewishvirtuallibrary.org', 'www.jcpa.org', 'ohelleah.org', 'jcckobe.org', 'www.jewishvirtuallibrary.org', 'www.kahaljoseph.org', 'dbs.bh.org', 'dbs.bh.org', 'jewishvirtuallibrary.org', 'www.jstor.org', 'www.jewishvirtuallibrary.org', 'www.jcpa.org', 'jewishvirtuallibrary.org', ['modern asian studies'], ['shofar'], ['proceedings of the american academy for jewish research']]",2206118,Allow all users (no expiry set),57387,10 July 2005,TShilo12 ,847,0,2005-07-10,2005-07,2005
560,560,North Malabar,https://en.wikipedia.org/wiki/North_Malabar,111,0,[],[],2,7,0,26,0,0,76,0.018018018018018018,0.06306306306306306,0.23423423423423423,0.0,0.0,0.08108108108108109,0,"['lsi.gov', 'censusindia.gov', 'lsi.gov', 'mahe.gov', 'lsi.gov', 'www.censusindia.gov', 'censusindia.gov', 'books.google.com', 'www.facebook.com', 'books.google.com', 'www.facesplacesandplates.com', 'books.google.com', 'ananthapuri.com', 'www.thehindu.com', 'www.thehindu.com', 'www.bbc.com', 'www.thehindu.com', 'recipesimply4u.blogspot.com', 'books.google.com', 'books.google.com', 'www.arabnews.com', 'books.google.com', 'deccanchronicle.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thetakeiteasychef.com', 'dcbookstore.com', 'books.google.com', 'books.google.com', 'www.legalserviceindia.com', 'www.deccanherald.com', 'www.cartage.org', 'krpcds.org']",22603905,Allow all users (no expiry set),82773,28 April 2009,Prakashkpc ,791,0,2009-04-28,2009-04,2009
561,561,Recife,https://en.wikipedia.org/wiki/Recife,108,0,[],[],16,32,0,48,0,0,13,0.14814814814814814,0.2962962962962963,0.4444444444444444,0.0,0.0,0.4444444444444444,0,"['www.inmet.gov', 'ftp.ibge.gov', 'www2.recife.pe.gov', 'cidades.ibge.gov', 'www.sidra.ibge.gov', 'www.portais.pe.gov', 'www.inmet.gov', 'www.inmet.gov', 'cidades.ibge.gov', 'geoftp.ibge.gov', 'www.recife.pe.gov', 'www.fundaj.gov', 'saladeimprensa.ibge.gov', 'www.inmet.gov', 'www.censo2010.ibge.gov', 'recife.pe.gov', 'www.cbtu.gov', 'www.inmet.gov', 'www.condepefidem.pe.gov', 'www.inmet.gov', 'www.censo2010.ibge.gov', 'www.cidades.ibge.gov', 'www.recife.pe.gov', 'www.inmet.gov', 'www.inmet.gov', 'www.inmet.gov', 'www.detran.pe.gov', 'basilio.fundaj.gov', 'www.recife.pe.gov', 'www.inmet.gov', 'basilio.fundaj.gov', 'www.inmet.gov', 'www.geographia.com', 'enotes.com', 'noticias.uol.com', 'www.brazil4you.com', 'www.cityknown.com', 'www.bbc.com', 'www.architecturaldigest.com', 'www.diariodepernambuco.com', 'www3.folhape.com', 'super.abril.com', 'blogs.diariodepernambuco.com', 'www2.uol.com', 'www2.uol.com', 'guiadolitoral.uol.com', 'congressoemfoco.uol.com', 'communis.com', 'www.aondefica.com', 'g1.globo.com', 'jc.uol.com', 'gwm2pub1.fishy.com', 'riomarrecife.com', 'oriettagggo.us.splinder.com', 'www.businessweek.com', 'www.caribbeannewsdigital.com', 'www.plazacasaforte.com', 'www.sharkattackdata.com', 'www.pernambuco.com', 'www.history.com', 'shoppingtacaruna.com', 'enotes.com', 'www.recifehotels.brazilhotels.4k.com', 'www.nassauturismo.com', 'www.projetocriancafelizbrasil.com', 'moovitapp.com', 'noticias.terra.com', 'viajandocomvoce.com', 'jconline.ne10.uol.com', 'www.geographia.com', 'oglobo.globo.com', 'www.recife.com', 'www.cine-pe.com', 'moovitapp.com', 'othersiderainbow.blogspot.com', 'blogs.diariodepernambuco.com', 'alljewishlinks.com', 'g1.globo.com', 'www.pe-az.com', 'www.diariodepernambuco.com', 'www.seguridadjusticiaypaz.org', 'ich.unesco.org', 'pt.wikipedia.org', 'www.globalvoicesonline.org', 'www.atlasbrasil.org', 'ich.unesco.org', 'whc.unesco.org', 'www.catholic-hierarchy.org', 'whc.unesco.org', 'www.portodigital.org', 'globalvoicesonline.org', 'www.redeandibrasil.org', 'creativecommons.org', 'www.blog.educacaoeparticipacao.org', 'ww2.panaftosa.org', 'www.cdsid.org']",65670,Allow all users (no expiry set),109032,29 July 2002,200.199.23.105 ,3335,5,2002-07-29,2002-07,2002
562,562,Afro-Dominicans,https://en.wikipedia.org/wiki/Afro-Dominicans,53,2,"['10.1080/00064246.2015.1060690', '10.5354/0719-4862.2018.50855', None, None, None, None]","[['black scholar '], ['meridional']]",7,3,0,21,0,0,20,0.1320754716981132,0.05660377358490566,0.39622641509433965,0.03773584905660377,0.0,0.22641509433962265,2,"['www.cia.gov', 'www.cia.gov', 'www.agn.gov', 'www.listindiario.com', 'www.nbcnews.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.listindiario.com', 'theroot.com', 'horacero.com', 'www.jmarcano.com', 'www.colonialzone-dr.com', 'ahorasecreto.blogspot.com', 'historiadominicana.com', 'diariolibre.com', 'www.buenastareas.com', 'books.google.com', 'www.listindiario.com', 'mindspring.com', 'www.caribbeannetnews.com', 'www.scribd.com', 'www.smithsonianmag.com', 'www.washingtonpost.com', 'innovation.org', 'www.oas.org', 'firstblacks.org', 'firstblacks.org', 'www.worldcat.org', 'antislavery.org', 'www.refworld.org', ['black scholar '], ['meridional']]",3106851,Allow all users (no expiry set),56887,8 November 2005,65.9.52.19 ,1302,5,2005-11-08,2005-11,2005
563,563,Sri Muktsar Sahib,https://en.wikipedia.org/wiki/Sri_Muktsar_Sahib,44,0,[],[],1,6,0,27,0,0,10,0.022727272727272728,0.13636363636363635,0.6136363636363636,0.0,0.0,0.1590909090909091,0,"['www.censusindia.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'censusindia.gov', 'agripb.gov', 'punjabjudiciary.gov', 'www.business-standard.com', 'www.mykhel.com', 'www.tribuneindia.com', 'www.urdupoint.com', 'punjabizm.com', 'www.historicalgurudwaras.com', 'www.dayandnightnews.com', 'www.worldgurudwaras.com', 'www.srimuktsarsahibonline.com', 'tribuneindia.com', 'www.worldgurudwaras.com', 'www.ndtv.com', 'yespunjab.com', 'www.hindustantimes.com', 'timesofindia.indiatimes.com', 'archive.indianexpress.com', 'archive.indianexpress.com', 'www.hoparoundindia.com', 'www.hindustantimes.com', 'www.sikhnugget.com', 'www.hindustantimes.com', 'mapsofindia.com', 'maplandia.com', 'www.highereducationinindia.com', 'www.worldgurudwaras.com', 'cricbuzz.com', 'www.hoparoundindia.com', 'oar.icrisat.org']",5802634,Allow all users (no expiry set),41306,2 July 2006,Ganeshbot ,663,0,2006-07-02,2006-07,2006
564,564,Christmas traditions,https://en.wikipedia.org/wiki/Christmas_traditions,69,0,[],[],7,1,0,20,0,0,42,0.10144927536231885,0.014492753623188406,0.2898550724637681,0.0,0.0,0.11594202898550725,0,"['schoolnet.gov', 'gbod-assets.s3.amazonaws.com', 'citybeat.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.italymagazine.com', 'www.christianitytoday.com', 'books.google.com', 'snopes.com', 'skiathosbooks.com', 'www.christmasarchives.com', 'books.google.com', 'www.etymonline.com', 'simplytreasures.com', 'books.google.com', 'books.google.com', 'www.fashion-era.com', 'www.boston.com', 'books.google.com', 'books.google.com', 'mistletoe.org', 'wayback.archive-it.org', 'www.catholicculture.org', 'www.npr.org', 'carnegiemnh.org', 'livius.org', 'www.saintnicholassociety.org']",62533138,Allow all users (no expiry set),52855,8 December 2019,Crumpled Fire ,57,0,2019-12-08,2019-12,2019
565,565,Kodava people,https://en.wikipedia.org/wiki/Kodava_people,90,0,[],[],0,3,0,54,0,0,33,0.0,0.03333333333333333,0.6,0.0,0.0,0.03333333333333333,0,"['pib.gov', 'censusindia.gov', 'censusindia.gov', 'books.google.com', 'www.deccanherald.com', 'www.hinduonnet.com', 'www.deccanherald.com', 'www.deccanherald.com', 'books.google.com', 'www.dnaindia.com', 'www.livemint.com', 'www.deccanherald.com', 'starofmysore.com', 'www.thehindu.com', 'www.coorgtourisminfo.com', 'wap.business-standard.com', 'www.deccanherald.com', 'www.thehindu.com', 'english.mathrubhumi.com', 'www.thehindu.com', 'www.coorg.com', 'www.newindianexpress.com', 'www.deccanherald.com', 'www.hinduonnet.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'www.evolveback.com', 'www.hindustantimes.com', 'm.economictimes.com', 'www.hinduonnet.com', 'www.thenewsminute.com', 'www.hinduonnet.com', 'www.deccanherald.com', 'www.deccanherald.com', 'motoxindia.com', 'www.hindu.com', 'books.google.com', 'www.newsncr.com', 'www.thehindu.com', 'www.thehindu.com', 'www.deccanherald.com', 'books.google.com', 'books.google.com', 'karnataka.com', 'www.deccanherald.com', 'www.thehindu.com', 'languageindia.com', 'www.hinduonnet.com', '0.gravatar.com', 'www.hindustantimes.com', 'www.britannica.com', 'books.google.com', 'www.hinduonnet.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.thehindu.com']",1456243,Allow all users (no expiry set),75261,1 February 2005,203.195.196.66 ,1687,5,2005-02-01,2005-02,2005
566,566,Homs,https://en.wikipedia.org/wiki/Homs,182,2,"['org/10.1017/cbo9780511676413', '10.3406/syria.1952.4788', None, None, None, None]","[['cambridge university press'], [' syria ']]",12,1,0,49,0,0,118,0.06593406593406594,0.005494505494505495,0.2692307692307692,0.01098901098901099,0.0,0.08241758241758242,2,"['www.dgam.gov', 'parsine.com', 'books.google.com', 'books.google.com', 'www.kadmusarts.com', 'en.oxforddictionaries.com', 'agha-syria.com', 'books.google.com', 'www.en.syria-scope.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'portalbelohorizonte.com', 'books.google.com', 'almaany.com', 'books.google.com', 'books.google.com', 'books.google.com', 'reference.allrefer.com', 'books.google.com', 'books.google.com', 'www.homsonline.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.weltfussballarchiv.com', 'www.collinsdictionary.com', 'www.cortasco.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.liilas.com', 'books.google.com', 'www.discover-syria.com', 'www.homsonline.com', 'www.bbc.com', 'books.google.com', 'www.kadmusarts.com', 'glosbe.com', 'worldpopulationreview.com', 'books.google.com', 'britannica.com', 'www.syriaphotoguide.com', 'www.weltfussballarchiv.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.newadvent.org', 'weekly.ahram.org', 'www.homscitycouncil.org', 'www.alnap.org', 'www.homscitycouncil.org', 'journals.openedition.org', 'www.cbssyr.org', 'www.homscitycouncil.org', 'www.homschamber.org', 'www.homscitycouncil.org', 'syriadirect.org', 'www.livius.org', ['cambridge university press'], [' syria ']]",77533,Allow all users (no expiry set),102589,29 August 2002,XJaM ,1827,9,2002-08-29,2002-08,2002
567,567,Entrevaux,https://en.wikipedia.org/wiki/Entrevaux,2,0,[],[],0,0,0,0,0,0,2,0.0,0.0,0.0,0.0,0.0,0.0,0,[],3124755,Allow all users (no expiry set),7033,10 November 2005,Olivier ,113,0,2005-11-10,2005-11,2005
568,568,Mantua,https://en.wikipedia.org/wiki/Mantua,11,0,[],[],0,1,0,2,0,0,8,0.0,0.09090909090909091,0.18181818181818182,0.0,0.0,0.09090909090909091,0,"['comune.mantova.gov', 'thewest.com', 'www.encyclopedia.com']",50187,Allow all users (no expiry set),30414,23 April 2002,65.30.64.186 ,818,1,2002-04-23,2002-04,2002
569,569,Culture of Afghanistan,https://en.wikipedia.org/wiki/Culture_of_Afghanistan,44,1,"['10.2307/521889', None, None]",[[' alif']],4,4,0,27,0,0,8,0.09090909090909091,0.09090909090909091,0.6136363636363636,0.022727272727272728,0.0,0.20454545454545456,1,"['photos.state.gov', 'lcweb2.loc.gov', 'www.cia.gov', 'afghanistan.usaid.gov', 'www.afghan-web.com', 'afghanmagazine.com', 'www.afghan-web.com', 'www.euppublishing.com', 'www.afghanproverbs.com', 'www.youtube.com', 'www.britannica.com', 'waronterrornews.typepad.com', 'www.foxnews.com', 'www.afghan-web.com', 'afghanmagazine.com', 'www.youtube.com', 'books.google.com', 'www.thehindubusinessline.com', 'about-afghanistan.squarespace.com', 'www.csmonitor.com', 'amp.theaustralian.com', 'www.tolonews.com', 'www.afghanistan-culture.com', 'www.bbc.com', 'www.awn.com', 'www.afghanproverbs.com', 'www.afghanproverbs.com', 'edition.cnn.com', 'www.afghanproverbs.com', 'www.pajhwok.com', 'www.sfgate.com', 'cp.settlement.org', 'www.pewforum.org', 'us.skateistan.org', 'newint.org', [' alif']]",1929224,Allow all users (no expiry set),33708,23 May 2005,Falphin ,1756,4,2005-05-23,2005-05,2005
570,570,Vlachs of Serbia,https://en.wikipedia.org/wiki/Vlachs_of_Serbia,67,0,[],[],10,5,0,7,0,0,45,0.14925373134328357,0.07462686567164178,0.1044776119402985,0.0,0.0,0.22388059701492538,0,"['webrzs.stat.gov', 'webrzs.stat.gov', 'webrzs.stat.gov', 'webrzs.stat.gov', 'webrzs.stat.gov', 'www.dw.com', 'www.glas-zajecara.com', 'www.britannica.com', 'books.google.com', 'www.vdss-petrovac.com', 'www.zajednicavlahasrbije.com', 'www.vdss-petrovac.com', 'www.timoc.org', 'fer.org', 'eparhija-timocka.org', 'www.isac-fund.org', 'www.arhivja.org', 'www.eparhijabihackopetrovacka.org', 'eparhija-timocka.org', 'fer.org', 'www.gergina.org', 'fer.org']",2888901,Allow all users (no expiry set),35663,12 October 2005,Ronline ,1234,7,2005-10-12,2005-10,2005
571,571,"Van, Turkey","https://en.wikipedia.org/wiki/Van,_Turkey",60,7,"['10.23976/smep.2014008', '10.1016/j.cscm.2015.10.001', '10.1080/13530199608705620', '10.1017/s0075435800066946', '10.1086/ahr/90.1.191-a', None, None, None, None, None, None, None, None, None, None]","[['singapore middle east papers'], ['case studies in construction materials'], ['british journal of middle eastern studies', 'taylor '], ['journal of roman studies'], ['the american historical review']]",5,2,0,14,0,0,32,0.08333333333333333,0.03333333333333333,0.23333333333333334,0.11666666666666667,0.0,0.23333333333333334,5,"['report.tuik.gov', 'www.mgm.gov', 'books.google.com', 'www.bbc.com', 'vanhavadis.com', 'vanhavadis.com', 'books.google.com', 'www.sophenearmeniaca.com', 'rbedrosian.com', 'www.hurriyetdailynews.com', 'www.armenian-history.com', 'edition.cnn.com', 'www.cnn.com', 'books.google.com', 'www.vangazetesi.com', 'www.sophenearmeniaca.com', 'www.metmuseum.org', 'books.openedition.org', 'www.iranicaonline.org', 'www.hrw.org', 'www.tesev.org', ['singapore middle east papers'], ['case studies in construction materials'], ['british journal of middle eastern studies', 'taylor '], ['journal of roman studies'], ['the american historical review']]",63685,Allow all users (no expiry set),43764,23 July 2002,imported>99.81,1772,8,2002-07-23,2002-07,2002
572,572,Valladolid,https://en.wikipedia.org/wiki/Valladolid,42,2,"['10.3989/estgeogr.201403', '10.5209/rev_docu.2016.v14.52898', None, None, None, None]","[['[[consejo superior de investigaciones científicas', 'estudios geográficos'], ['documenta ', '[[complutense university of madrid']]",2,0,0,7,0,0,31,0.047619047619047616,0.0,0.16666666666666666,0.047619047619047616,0.0,0.09523809523809523,2,"['rsssf.com', 'www.xlsemanal.com', 'www.lavanguardia.com', 'elpais.com', 'www.romanicodigital.com', 'www.tribunasalamanca.com', 'www.lavanguardia.com', 'lfcyl.org', 'books.openedition.org', ['[[consejo superior de investigaciones científicas', 'estudios geográficos'], ['documenta ', '[[complutense university of madrid']]",69311,Allow all users (no expiry set),57491,8 August 2002,207.253.140.103 ,1305,6,2002-08-08,2002-08,2002
573,573,South Malabar,https://en.wikipedia.org/wiki/South_Malabar,219,3,"['10.2307/2690896', '10.1086/356288', None, None, None, None]","[['mathematics magazine '], ['isis ']]",23,24,0,103,0,0,66,0.1050228310502283,0.1095890410958904,0.4703196347031963,0.0136986301369863,0.0,0.228310502283105,2,"['sametham.kite.kerala.gov', 'spb.kerala.gov', 'nielit.gov', 'industry.kerala.gov', 'lsi.gov', 'sametham.kite.kerala.gov', 'lsi.gov', 'www.mlp.kerala.gov', 'censusindia.gov', 'www.prd.kerala.gov', 'sametham.kite.kerala.gov', 'censusindia.gov', 'sametham.kite.kerala.gov', 'dmg.kerala.gov', 'lsi.gov', 'sametham.kite.kerala.gov', 'censusindia.gov', 'sametham.kite.kerala.gov', 'spb.kerala.gov', 'sametham.kite.kerala.gov', 'ecostat.kerala.gov', 'www.kkd.kerala.gov', 'sametham.kite.kerala.gov', 'www.igcar.gov', 'thehindu.com', 'facesplacesandplates.com', 'www.deccanchronicle.com', 'gulfnews.com', 'www.business-standard.com', 'www.thehindu.com', 'mighil.com', 'english.forbesmiddleeast.com', 'www.newindianexpress.com', 'books.google.com', 'webindia123.com', 'www.thehindu.com', 'www.thehindubusinessline.com', 'www.thehindu.com', 'english.manoramaonline.com', 'articles.timesofindia.indiatimes.com', 'articles.timesofindia.indiatimes.com', 'cricketarchive.com', 'www.thehindu.com', 'www.thehindu.com', 'www.newindianexpress.com', 'www.thehindu.com', 'www.hindu.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'rediff.com', 'thehindu.com', 'kozhikode.cyberparktoday.com', 'www.thehindubusinessline.com', 'nilamburnews.com', 'books.google.com', 'manoramaonline.com', 'www.mathrubhumi.com', 'www.manoramaonline.com', 'www.thehindu.com', 'www.thehindu.com', 'www.mathrubhumi.com', 'hellobahrain.com', 'www.hindu.com', 'thehindu.com', 'www.thehindu.com', 'oonmanorama.com', 'articles.timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'india.com', 'www.asianage.com', 'english.mathrubhumi.com', 'thehindu.com', 'www.cookawesome.com', 'www.calicutpressclub.com', 'www.thehindu.com', 'post.artoflegendindia.com', 'timesofindia.indiatimes.com', 'www.variety.com', 'www.mathrubhumi.com', 'www.thehindu.com', 'www.deccanchronicle.com', 'puzhakal0.tripod.com', 'timesofindia.indiatimes.com', 'www.hindu.com', 'espncricinfo.com', 'www.yatra.com', 'www.thehindu.com', 'imsmagic.com', 'www.thehindu.com', 'english.mathrubhumi.com', 'www.deccanchronicle.com', 'timesofindia.indiatimes.com', 'onmanorama.com', 'books.google.com', 'kozhikode.com', 'www.mathrubhumi.com', 'timesofindia.indiatimes.com', 'www.newindianexpress.com', 'www.newindianexpress.com', 'www.vccircle.com', 'articles.timesofindia.indiatimes.com', 'thiraseela.com', 'www.hindu.com', 'dcbookstore.com', 'businesswireindia.com', 'books.google.com', 'timesofindia.indiatimes.com', 'www.mapsofindia.com', 'www.thehindu.com', 'timesofindia.indiatimes.com', 'aryavaidyasala.com', 'www.arabnews.com', 'timesofindia.indiatimes.com', 'keralartc.com', 'www.thehindu.com', 'www.thehindu.com', 'www.ethnologue.com', 'books.google.com', 'epaper.malayalamvaarika.com', 'www.hindu.com', 'www.deccanchronicle.com', 'www.deccanherald.com', 'nwitimes.com', 'www.thehindu.com', 'diehardindian.com', 'www.hindu.com', 'nativeplanet.com', 'www.cartage.org', 'keralatourism.org', 'keralatourism.org', 'www.birdlife.org', 'keralatourism.org', 'keralasahityaakademi.org', 'keralatourism.org', 'keralatourism.org', 'keralatourism.org', 'malappuramtourism.org', 'keralaassembly.org', 'cmgmusiccollege.org', 'tyagaraja-aradhana-calicut.org', 'malappuramtourism.org', 'keralatourism.org', 'keralatourism.org', 'www.nhai.org', 'keralatourism.org', 'keralatourism.org', 'palakkadtourism.org', 'cyberparkkerala.org', 'www.keralatourism.org', 'keralatourism.org', ['mathematics magazine '], ['isis ']]",64652632,Allow all users (no expiry set),165759,26 July 2020,Kambliyil ,220,0,2020-07-26,2020-07,2020
574,574,Northeast China,https://en.wikipedia.org/wiki/Northeast_China,22,0,[],[],6,1,0,10,0,0,5,0.2727272727272727,0.045454545454545456,0.45454545454545453,0.0,0.0,0.3181818181818182,0,"['www.gov', 'andrewbatson.com', 'books.google.com', 'thediplomat.com', 'www.forbes.com', 'www.scmp.com', 'www.theatlantic.com', 'www.scmp.com', 'english.caixin.com', 'books.google.com', 'books.google.com', 'www.jstor.org', 'www.jstor.org', 'www.jstor.org', 'www.jstor.org', 'www.jstor.org', 'www.jstor.org']",788662,Allow all users (no expiry set),24432,6 July 2004,Ran ,586,5,2004-07-06,2004-07,2004
575,575,Culture of Egypt,https://en.wikipedia.org/wiki/Culture_of_Egypt,13,0,[],[],1,1,0,6,0,0,5,0.07692307692307693,0.07692307692307693,0.46153846153846156,0.0,0.0,0.15384615384615385,0,"['www.sis.gov', 'books.google.com', 'ukhotmovies.com', 'www.harvardmagazine.com', 'www.dawn.com', 'archive.fiba.com', 'archive.fiba.com', 'www.globalcitizen.org']",51218,Allow all users (no expiry set),32770,3 May 2002,Eclecticology ,1921,0,2002-05-03,2002-05,2002
576,576,Kavala,https://en.wikipedia.org/wiki/Kavala,30,0,[],[],2,0,0,6,0,0,22,0.06666666666666667,0.0,0.2,0.0,0.0,0.06666666666666667,0,"['www.kavala-airshow.com', 'www.kavala-cosmopolis.com', 'www.sistercities-durham.com', 'www.egnatia-aviation.com', 'gradgradiska.com', 'www.railjournal.com', 'www.ilak.org', 'www.mohamed-ali.org']",234317,Allow all users (no expiry set),44464,26 May 2003,217.155.80.220 ,1040,5,2003-05-26,2003-05,2003
577,577,Dodecanese,https://en.wikipedia.org/wiki/Dodecanese,21,2,"['10.1080/09592299308405886', '10.12681/eoaesperia.78', None, None, None, None]","[['diplomacy and statecraft '], [' ἑῶα καὶ ἑσπέρια ']]",1,1,0,5,0,0,12,0.047619047619047616,0.047619047619047616,0.23809523809523808,0.09523809523809523,0.0,0.19047619047619047,2,"['www.mfa.gov', 'www.sabah.com', 'books.google.com', 'www.johnhearfield.com', 'ng3k.com', 'books.google.com', 'www.eoearth.org', ['diplomacy and statecraft '], [' ἑῶα καὶ ἑσπέρια ']]",302628,Allow all users (no expiry set),34215,22 August 2003,195.242.150.176 ,633,0,2003-08-22,2003-08,2003
578,578,Northern Norway,https://en.wikipedia.org/wiki/Northern_Norway,37,1,"['10.1016/j.meatsci.2009.08.008', '20416633', None]",[['meat science ']],1,0,0,5,0,0,30,0.02702702702702703,0.0,0.13513513513513514,0.02702702702702703,0.0,0.05405405405405406,1,"['thebarentsobserver.com', 'www.newscientist.com', 'issuu.com', 'pickyourtrail.com', 'boknafisk.com', 'www.eu-interact.org', ['meat science ']]",1433683,Allow all users (no expiry set),61498,26 January 2005,Egil ,617,1,2005-01-26,2005-01,2005
579,579,Vendée,https://en.wikipedia.org/wiki/Vend%C3%A9e,11,0,[],[],0,0,0,2,0,0,9,0.0,0.0,0.18181818181818182,0.0,0.0,0.0,0,"['www.mareuiltourisme.com', 'books.google.com']",88951,Allow all users (no expiry set),22575,21 September 2002,209.105.200.23 ,504,0,2002-09-21,2002-09,2002
580,580,Jämtland,https://en.wikipedia.org/wiki/J%C3%A4mtland,38,0,[],[],2,0,0,4,0,0,32,0.05263157894736842,0.0,0.10526315789473684,0.0,0.0,0.05263157894736842,0,"['regionfakta.com', 'www.noside.com', 'www.jamtli.com', 'scotsman.com', 'jamtamot.org', 'www.verdal.historielag.org']",190814,Allow all users (no expiry set),81129,2 March 2003,Mic ,583,0,2003-03-02,2003-03,2003
581,581,Isleños (Louisiana),https://en.wikipedia.org/wiki/Isle%C3%B1os_(Louisiana),30,2,"['10.2307/2595192', '10.2307/335051', None, None, None, None]","[['the economic history review', 'wiley on behalf of the economic history society'], ['hispania']]",6,1,0,9,0,0,12,0.2,0.03333333333333333,0.3,0.06666666666666667,0.0,0.3,2,"['www.census.gov', 'www.theadvocate.com', 'www.wafb.com', 'nola.verylocal.com', 'www.google.com', 'www.newspapers.com', 'books.google.com', 'www.miamiherald.com', 'www.newspapers.com', 'www.nbcnews.com', 'www.canaryislanders.org', 'www.mackseysymposium.org', 'www.losislenos.org', 'projects.propublica.org', 'www.canaryislanders.org', 'www.losislenos.org', ['the economic history review', 'wiley on behalf of the economic history society'], ['hispania']]",45402537,Allow all users (no expiry set),41833,14 February 2015,Isinbill ,415,0,2015-02-14,2015-02,2015
582,582,Thalassery,https://en.wikipedia.org/wiki/Thalassery,54,1,"['10.2307/3516674', None, None]",[['social scientist ']],6,6,0,24,0,0,17,0.1111111111111111,0.1111111111111111,0.4444444444444444,0.018518518518518517,0.0,0.24074074074074073,1,"['prd.kerala.gov', 'mahe.gov', 'www.kerala.gov', 'censusindia.gov', 'india-wris.nrsc.gov', 'www.keralapwd.gov', 'hindu.com', 'articles.timesofindia.indiatimes.com', 'www.thehindu.com', 'www.spiceography.com', 'www.theyyamcalendar.com', 'articles.economictimes.indiatimes.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'hindustankalari.com', 'articles.timesofindia.indiatimes.com', 'www.mysingaporekitchen.com', 'www.kannurtourism.com', 'www.newindianexpress.com', 'www.hindu.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.worldweatheronline.com', 'www.thehindu.com', 'www.thehindu.com', 'www.keralacricketonline.com', 'epaper.newindianexpress.com', 'www.thehindu.com', 'gulfnews.com', 'www.thehindu.com', 'www.keralatourism.org', 'www.indiaenvironmentportal.org', 'www.kannurairport.org', 'www.keralatourism.org', 'www.keralatourism.org', 'en.climate-data.org', ['social scientist ']]",1235269,Allow all users (no expiry set),43003,2 December 2004,64.26.228.77 ,2586,14,2004-12-02,2004-12,2004
583,583,Gümüşhane,https://en.wikipedia.org/wiki/G%C3%BCm%C3%BC%C5%9Fhane,18,0,[],[],1,3,0,8,0,0,6,0.05555555555555555,0.16666666666666666,0.4444444444444444,0.0,0.0,0.2222222222222222,0,"['www.kulturturizm.gov', 'www.mgm.gov', 'report.tuik.gov', 'www.karalahana.com', 'karalahana.com', 'www.statoids.com', 'www.visiontours.com', 'www.fallingrain.com', 'www.karalahana.com', 'books.google.com', 'karalahana.com', 'www.wdl.org']",2581973,Allow all users (no expiry set),24264,31 August 2005,Macukali ,378,0,2005-08-31,2005-08,2005
584,584,Goan Catholics,https://en.wikipedia.org/wiki/Goan_Catholics,216,0,[],[],11,4,0,115,0,0,87,0.05092592592592592,0.018518518518518517,0.5324074074074074,0.0,0.0,0.06944444444444445,0,"['www.india.gov', 'www.india.gov', 'www.censusindia.gov', 'www.india.gov', 'm.timesofindia.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'content-www.cricinfo.com', 'www.daijiworld.com', 'books.google.com', 'hillmanwonders.com', 'm.timesofindia.com', 'books.google.com', 'm.timesofindia.com', 'www.hinduonnet.com', 'economictimes.indiatimes.com', 'books.google.com', 'www.daijiworld.com', 'www.hinduonnet.com', 'www.daijiworld.com', 'www.firstpost.com', 'books.google.com', 'books.google.com', 'www.hindu.com', 'books.google.com', 'www.konkanisongbook.com', 'books.google.com', 'books.google.com', 'books.google.com', 'indianfootball.com', 'www.navhindtimes.com', 'groups.yahoo.com', 'www.hindu.com', 'books.google.com', 'indianexpress.com', 'books.google.com', 'books.google.com', 'www.merinews.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.ethnologue.com', 'books.google.com', 'books.google.com', 'www.patriciarozario.com', 'www.hinduonnet.com', 'books.google.com', 'books.google.com', 'www.goansinoman.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.hindu.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.deccanherald.com', 'www.navhindtimes.com', 'goacom.com', 'www.india-today.com', 'www.flickr.com', 'books.google.com', 'goacom.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'books.google.com', 'www.daijiworld.com', 'www.goatoronto.com', 'books.google.com', 'books.google.com', 'www.dawn.com', 'books.google.com', 'm.timesofindia.com', 'books.google.com', 'm.timesofindia.com', 'www.dnaindia.com', 'keithvaz.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.goatoronto.com', 'books.google.com', 'books.google.com', 'articles.timesofindia.indiatimes.com', 'gulfnews.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.hindu.com', 'www.mail-archive.com', 'books.google.com', 'books.google.com', 'books.google.com', 'timesofindia.indiatimes.com', 'books.google.com', 'books.google.com', 'www.tehelka.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.goacom.com', 'the-aiff.com', 'books.google.com', 'books.google.com', 'abbefaria.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.goanvoice.org', 'www.portcities.org', 'infochangeindia.org', 'www.goanvoice.org', 'www.portcities.org', 'www.goatourism.org', 'www.ylgs.org', 'www.archbom.org', 'lists.goanet.org', 'www.goakonkaniakademi.org', 'americancatholic.org']",5931351,Allow all users (no expiry set),89261,12 July 2006,Hornplease ,5481,2,2006-07-12,2006-07,2006
585,585,Afro–Puerto Ricans,https://en.wikipedia.org/wiki/Afro%E2%80%93Puerto_Ricans,137,7,"['10.1371/journal.pone.0016513', '10.2307/2571712', '10.1353/hcs.2007.0017', '10.1177/000312240707200604', '10.14452/mr-055-10-2004-03_1', '10.2307/2574293', '21304981', None, None, None, None, None, '3031579', None, None, None, None, None]","[['plos one '], ['social forces '], ['arizona journal of hispanic cultural studies '], ['american sociological review '], ['monthly review '], ['social forces ']]",12,9,0,71,0,0,38,0.08759124087591241,0.06569343065693431,0.5182481751824818,0.051094890510948905,0.0,0.20437956204379562,6,"['2010.census.gov', 'loc.gov', 'www.census.gov', 'www.loc.gov', 'www.census.gov', 'census.gov', 'factfinder.census.gov', 'www.loc.gov', 'cia.gov', 'caribbeanbusinesspr.com', 'books.google.com', 'hispanicallyspeakingnews.com', 'angelfire.com', 'cwo.com', 'allaboutjazz.com', 'proyectosalonhogar.com', 'huffingtonpost.com', 'latino.foxnews.com', 'tracingafricanroots.wordpress.com', 'www.fortunecity.com', 'tracingafricanroots.wordpress.com', 'usatoday.com', 'shagtown.com', 'fortunecity.com', 'espn.go.com', 'www.ibhof.com', 'encantada2006.blogspot.com', 'vocero.com', 'www.fortunecity.com', 'blackvoicenews.com', 'triplov.com', 'ipoaa.com', 'hipsonfire.com', 'boston.com', 'encantada2006.blogspot.com', 'cubacreme.com', 'zonai.com', 'caribbeantrading.com', 'www.cbsnews.com', 'stewartsynopsis.com', 'angelfire.com', 'www.nlbpa.com', 'triplov.com', 'elliesbookz.wordpress.com', 'kwekudee-tripdownmemorylane.blogspot.com', 'rain-people.com', 'tracingafricanroots.wordpress.com', 'indexarticles.com', 'www.newspapers.com', 'nylatinojournal.com', 'fullbooks.com', 'books.google.com', 'linktopr.com', 'preb.com', 'caribbeantrading.com', 'elliesbookz.wordpress.com', 'www.ipoaa.com', 'shagtown.com', 'repeatingislands.com', 'www.nydailynews.com', 'cwo.com', 'tracingafricanroots.wordpress.com', 'nativetimes.com', 'www.timboucher.com', 'kwekudee-tripdownmemorylane.blogspot.com', 'stewartsynopsis.com', 'www.rhythmweb.com', 'www.nydailynews.com', 'indexarticles.com', 'finalcall.com', 'tracingafricanroots.wordpress.com', 'proyectosalonhogar.com', 'www.musicofpuertorico.com', 'www.ew.com', 'ipoaa.com', 'sportsillustrated.cnn.com', 'www.seeingblack.com', 'xpertia.com', 'tracingafricanroots.wordpress.com', 'fortunecity.com', 'www.losplenerosdela21.org', 'www.npr.org', 'www.afropedea.org', 'www.puertorico-herald.org', 'firstblacks.org', 'latinousa.org', 'prpop.org', 'minorityrights.org', 'oecd.org', 'ensayistas.org', 'minorityrights.org', 'www.npr.org', ['plos one '], ['social forces '], ['arizona journal of hispanic cultural studies '], ['american sociological review '], ['monthly review '], ['social forces ']]",4517597,Allow all users (no expiry set),96849,26 March 2006,Marine 69-71 ,1459,28,2006-03-26,2006-03,2006
586,586,Tokat,https://en.wikipedia.org/wiki/Tokat,10,0,[],[],1,2,0,3,0,0,4,0.1,0.2,0.3,0.0,0.0,0.3,0,"['www.mgm.gov', 'www2.diyanet.gov', 'www.tokatgazetesi.com', 'www.huffingtonpost.com', 'pontosworld.com', 'www.jstor.org']",1337996,Allow all users (no expiry set),15898,28 December 2004,Llywrch ,344,0,2004-12-28,2004-12,2004
587,587,Syrian Jews,https://en.wikipedia.org/wiki/Syrian_Jews,46,0,[],[],5,0,0,24,0,0,17,0.10869565217391304,0.0,0.5217391304347826,0.0,0.0,0.10869565217391304,0,"['www.cnn.com', 'www.youtube.com', 'ninemonthsinsyria.blogspot.com', 'www.youtube.com', 'www.nytimes.com', 'books.google.com', 'www.timesofisrael.com', 'www.israelfaxx.com', 'www.nytimes.com', 'www.jpost.com', 'www.nytimes.com', 'www.nytimes.com', 'www.vosizneias.com', 'www.nytimes.com', 'books.google.com', 'recipelink.com', 'www.shaar-binyamin.com', 'www.simpletoremember.com', 'wsj.com', 'www.al-monitor.com', 'www.jpost.com', 'jewishencyclopedia.com', 'www.simpletoremember.com', 'www.aleppojews.com', 'www.nli.org', 'digital.cjh.org', 'www.jewishvirtuallibrary.org', 'www.jewishvirtuallibrary.org', 'www.piyut.org']",5531820,Allow all users (no expiry set),57295,12 June 2006,Sirmylesnagopaleentheda ,2496,1,2006-06-12,2006-06,2006
588,588,Jewish culture,https://en.wikipedia.org/wiki/Jewish_culture,129,2,"['10.1353/ajh.2015.0023', '10.1038/187493a0', None, None, None, None]","[['american jewish history'], ['nature ']]",26,0,0,54,0,1,47,0.20155038759689922,0.0,0.4186046511627907,0.015503875968992248,0.0,0.21705426356589147,2,"['forward.com', 'www.nbcnews.com', 'www.jewishencyclopedia.com', 'articles.washingtonpost.com', 'www.thejc.com', 'www.timesofisrael.com', 'www.timesofisrael.com', 'jewishencyclopedia.com', 'www.geocities.com', 'www.toonopedia.com', 'britannica.com', 'www.myjewishlearning.com', 'gme.grolier.com', 'books.google.com', 'willeisner.com', 'judaism.com', 'www.jewishjournal.com', 'www.diningchicago.com', 'www.tcj.com', 'www.ynetnews.com', 'www.gulf-daily-news.com', 'myjewishlearning.com', 'myjewishlearning.com', 'www.playbill.com', 'books.google.com', 'find.galegroup.com', 'query.nytimes.com', 'books.google.com', 'www.forward.com', 'forward.com', 'jewishencyclopedia.com', 'ralphbakshi.com', 'books.google.com', 'www.talkinbroadway.com', 'www.bonappetit.com', 'www.jewish-theatre.com', 'gme.grolier.com', 'www.policonomics.com', 'www.bbc.com', 'www.shalomlife.com', 'momentmag.com', 'select.nytimes.com', 'www.haaretz.com', 'myjewishlearning.com', 'gme.grolier.com', 'www.jewish-theatre.com', 'www.nature.com', 'www.toonopedia.com', 'amazon.com', 'books.google.com', 'www.haaretz.com', 'myjewishlearning.com', 'www.jewishsf.com', 'leonardbernstein.com', 'www.imj.org', 'www.jewishvirtuallibrary.org', 'www.bje.org', 'jinfo.org', 'livius.org', 'www.hadassah.org', 'habima.org', 'jinfo.org', 'www.pbs.org', 'meitar.org', 'www.thejewishmuseum.org', 'jinfo.org', 'www.jinfo.org', 'www.jmi.org', 'www.jewishvirtuallibrary.org', 'www.jinfo.org', 'www.sciencemuseum.org', 'www.jstor.org', 'jewishvirtuallibrary.org', 'www.jcpa.org', 'www.ejpress.org', 'www.dnaftb.org', 'www.jinfo.org', 'www.cjh.org', 'jinfo.org', 'www.machar.org', ['american jewish history'], ['nature ']]",1262063,Allow all users (no expiry set),125792,10 December 2004,IZAK ,1908,3,2004-12-10,2004-12,2004
589,589,Sardinian people,https://en.wikipedia.org/wiki/Sardinian_people,264,14,"['10.1093/molbev/msx082', '10.1038/s41467-020-14523-6', '10.1038/ng.3368', '10.1038/sj.ejcn.1602596', '10.1371/journal.pone.0190169', '10.1038/s41559-020-1102-0', '10.1371/journal.pone.0043759', '10.1038/ng.3426', '10.1046/j.1468-1331.2002.00412.x', '10.1371/journal.pone.0091237', '10.1159/000109884', None, '28177087', '32094358', '26366554', '17228351', '29320542', '32094539', '22984441', '26506900', '12099914', '24651212', '8719044', None, '5400395', '7039977', '4627508', None, '5761892', '7080320', '3440425', None, None, '3961211', None, None]","[[' mol. biol. evol. '], ['nature', 'nature communications'], ['nature genetics '], ['eur j clin nutr '], [' plos one', 'pubmed central'], ['nature ecology and evolution '], ['plos one'], [' nat. genet. '], ['eur j neurol '], ['plos one '], ['neuroepidemiology '], ['nature ecology ']]",6,0,0,33,0,2,208,0.022727272727272728,0.0,0.125,0.05303030303030303,0.0,0.07575757575757576,12,"['books.google.com', 'www.sardegnasoprattutto.com', 'www.degruyter.com', 'genographic.nationalgeographic.com', 'www.bluezones.com', 'www.cell.com', 'eupedia.com', 'www.nature.com', 'www.mdpi.com', 'books.google.com', 'books.google.com', 'www.bluezones.com', 'www.sciencedaily.com', 'www.nature.com', 'www.msdmanuals.com', 'www.thelatinlibrary.com', 'www.nature.com', 'thebark.com', 'seosardinia.wordpress.com', 'www.nature.com', 'www.etymonline.com', 'www.ethnologue.com', 'www.nature.com', 'www.nature.com', 'seosardinia.wordpress.com', 'maxia-mail.doomby.com', 'www.encyclopedia.com', 'www.nature.com', 'www.nature.com', 'www.bluezones.com', 'www.lexico.com', 'www.ethnologue.com', 'static-content.springer.com', 'mbe.oxfordjournals.org', 'science.sciencemag.org', 'biorxiv.org', 'www.unesco.org', 'www.genetics.org', 'www.refworld.org', [' mol. biol. evol. '], ['nature', 'nature communications'], ['nature genetics '], ['eur j clin nutr '], [' plos one', 'pubmed central'], ['nature ecology and evolution '], ['plos one'], [' nat. genet. '], ['eur j neurol '], ['plos one '], ['neuroepidemiology '], ['nature ecology ']]",27644194,Allow all users (no expiry set),112168,8 June 2010,Xoil ,1555,2,2010-06-08,2010-06,2010
590,590,Salzwedel,https://en.wikipedia.org/wiki/Salzwedel,2,0,[],[],0,0,0,0,0,0,2,0.0,0.0,0.0,0.0,0.0,0.0,0,[],162235,Allow all users (no expiry set),11042,28 December 2002,212.59.62.132 ,173,0,2002-12-28,2002-12,2002
591,591,Acireale,https://en.wikipedia.org/wiki/Acireale,4,0,[],[],0,0,0,1,0,0,3,0.0,0.0,0.25,0.0,0.0,0.0,0,['www.com'],1547513,Allow all users (no expiry set),13241,26 February 2005,J heisenberg ,281,0,2005-02-26,2005-02,2005
592,592,List of English words of Italian origin,https://en.wikipedia.org/wiki/List_of_English_words_of_Italian_origin,32,0,[],[],1,0,0,23,0,0,8,0.03125,0.0,0.71875,0.0,0.0,0.03125,0,"['www.etymonline.com', 'www.etymonline.com', 'www.etymonline.com', 'www.etymonline.com', 'www.etymonline.com', 'www.etymonline.com', 'www.etymonline.com', 'www.etymonline.com', 'www.etymonline.com', 'www.etymonline.com', 'www.etymonline.com', 'www.etymonline.com', 'www.etymonline.com', 'www.etymonline.com', 'www.thelmagazine.com', 'www.etymonline.com', 'dictionary.reference.com', 'www.myetymology.com', 'www.etymonline.com', 'oxforddictionaries.com', 'www.etymonline.com', 'worldsoccer.com', 'www.etymonline.com', 'www.worldwidewords.org']",39432784,Allow all users (no expiry set),28268,20 May 2013,Grutness ,285,2,2013-05-20,2013-05,2013
593,593,History of the Jews in Thessaloniki,https://en.wikipedia.org/wiki/History_of_the_Jews_in_Thessaloniki,70,1,"['10.1093/hgs/14.2.165', None, None]",[['holocaust and genocide studies']],8,1,0,5,0,0,55,0.11428571428571428,0.014285714285714285,0.07142857142857142,0.014285714285714285,0.0,0.14285714285714285,1,"['www.state.gov', 'www.orbilat.com', 'www.routledge.com', 'www.orbilat.com', 'greece.greekreporter.com', 'greekreporter.com', 'dbs.bh.org', 'www.etzahaim.org', 'www.akadem.org', 'faktencheckhellas.org', 'fmh.org', 'www.ushmm.org', 'www.jta.org', 'hts.org', ['holocaust and genocide studies']]",14030921,Allow all users (no expiry set),79972,2 November 2007,Eliyak ,814,1,2007-11-02,2007-11,2007
594,594,Kastoria,https://en.wikipedia.org/wiki/Kastoria,36,0,[],[],4,0,0,10,0,0,22,0.1111111111111111,0.0,0.2777777777777778,0.0,0.0,0.1111111111111111,0,"['trezoros.com', 'books.google.com', 'www.nytimes.com', 'www.plovdivguide.com', 'www.nytimes.com', 'dictionary.oed.com', 'greekreporter.com', 'hauteacorn.com', 'greece.greekreporter.com', 'www.timesofisrael.com', 'jewishvirtuallibrary.org', 'www.ushmm.org', 'www.promacedonia.org', 'www.jstor.org']",302636,Allow all users (no expiry set),37503,22 August 2003,195.242.150.176 ,1081,6,2003-08-22,2003-08,2003
595,595,"Cáceres, Spain","https://en.wikipedia.org/wiki/C%C3%A1ceres,_Spain",22,1,"['10.1126/science.aap7778', '29472483', None]",[['science ']],3,0,0,4,0,1,13,0.13636363636363635,0.0,0.18181818181818182,0.045454545454545456,0.0,0.18181818181818182,1,"['www.elperiodicoextremadura.com', 'www.elperiodicoextremadura.com', 'www.irishfleadhcaceres.com', 'www.elperiodicoextremadura.com', 'ab.dip-caceres.org', 'www.turismocaceres.org', 'thesession.org', ['science ']]",143655,Allow all users (no expiry set),25401,3 November 2002,Montrealais ,441,0,2002-11-03,2002-11,2002
596,596,History of Indian influence on Southeast Asia,https://en.wikipedia.org/wiki/History_of_Indian_influence_on_Southeast_Asia,124,4,"['10.1038/s41598-018-22995-2', '10.7152/bippa.v30i0.9966', '10.1038/nature21696', '10.1179/014703783788755502', '29581431', None, '28277506', None, '5979964', None, None, None]","[['scientific reports'], ['bulletin of the indo-pacific prehistory association ', ' indo-pacific prehistory association '], ['nature'], [' ming studies ']]",5,4,0,29,0,0,82,0.04032258064516129,0.03225806451612903,0.23387096774193547,0.03225806451612903,0.0,0.10483870967741936,4,"['state.gov', 'www.nla.gov', 'eresources.nlb.gov', 'eresources.nlb.gov', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.cebu-online.com', 'www.southeastasianarchaeology.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.zambotoday.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.seaarchaeology.com', 'books.google.com', 'anaknabinalatongan.wixsite.com', 'books.google.com', 'books.google.com', 'www.silk-road.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.esamskriti.com', 'www.mathrubhumi.com', 'books.google.com', 'books.google.com', 'www.reninc.org', 'www.reninc.org', 'www.khmerstudies.org', 'www.pbs.org', 'www.oocities.org', ['scientific reports'], ['bulletin of the indo-pacific prehistory association ', ' indo-pacific prehistory association '], ['nature'], [' ming studies ']]",38028031,Allow all users (no expiry set),112536,26 December 2012,Irahulpandey ,339,4,2012-12-26,2012-12,2012
597,597,Piana degli Albanesi,https://en.wikipedia.org/wiki/Piana_degli_Albanesi,41,1,"['10.1093/pastj/gtq030', None, None]",[['past ']],2,0,0,4,0,0,34,0.04878048780487805,0.0,0.0975609756097561,0.024390243902439025,0.0,0.07317073170731707,1,"['books.google.com', 'www.com', 'booksandjournals.brillonline.com', 'books.google.com', 'gcatholic.org', 'www.balcanicaucaso.org', ['past ']]",5588157,Allow all users (no expiry set),52772,16 June 2006,Djalo24 ,738,1,2006-06-16,2006-06,2006
598,598,Syros,https://en.wikipedia.org/wiki/Syros,17,0,[],[],0,0,0,4,0,0,13,0.0,0.0,0.23529411764705882,0.0,0.0,0.0,0,"['www.turkcebilgi.com', 'greeka.com', 'books.google.com', 'www.economist.com']",276987,Allow all users (no expiry set),28052,25 July 2003,194.219.81.125 ,662,0,2003-07-25,2003-07,2003
599,599,Tabriz,https://en.wikipedia.org/wiki/Tabriz,134,5,"['10.1080/05786967.2007.11864720', '10.1080/713687484', '10.22034/gjesm.2018.04.02.007', None, None, None, None, None, None]","[['iran'], ['nationalities papers ', (' nationalities papers', ' papers', 'papers', 'v')], ['global journal of environmental science and management ']]",13,1,0,28,0,0,88,0.09701492537313433,0.007462686567164179,0.208955223880597,0.03731343283582089,0.0,0.1417910447761194,3,"['in.gov', 'brill.com', 'www.iotpe.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'asreazadi.com', 'www.encyclopaediaislamica.com', 'www.mehrnews.com', 'www.tavoosonline.com', 'articles.businessinsider.com', 'www.farsnews.com', 'farsnews.com', 'books.google.com', 'www.britannica.com', 'rsssf.com', 'books.google.com', 'books.google.com', 'www.farsnews.com', 'books.google.com', 'books.google.com', 'www.worldclimate.com', 'www.magiran.com', 'concise.britannica.com', 'books.google.com', 'www.farsnews.com', 'www.farsnews.com', 'electricpulp.com', 'www.iranicaonline.org', 'www.amar.org', 'amar.sci.org', 'realiran.org', 'sci.org', 'www.amar.org', 'sci.org', 'www.amar.org', 'www.prsir.org', 'tabrizcity.org', 'whc.unesco.org', 'wccapr.org', 'www.iranicaonline.org', ['iran'], ['nationalities papers ', (' nationalities papers', ' papers', 'papers', 'v')], ['global journal of environmental science and management ']]",439791,Allow all users (no expiry set),108723,23 January 2004,DigiBullet ,5646,4,2004-01-23,2004-01,2004
600,600,Niksar,https://en.wikipedia.org/wiki/Niksar,8,0,[],[],1,0,0,2,0,0,5,0.125,0.0,0.25,0.0,0.0,0.125,0,"['books.google.com', 'books.google.com', 'whc.unesco.org']",2760424,Allow all users (no expiry set),14433,25 September 2005,145.99.193.143 ,225,1,2005-09-25,2005-09,2005
601,601,"Bellagio, Lombardy","https://en.wikipedia.org/wiki/Bellagio,_Lombardy",29,0,[],[],3,0,0,2,0,0,24,0.10344827586206896,0.0,0.06896551724137931,0.0,0.0,0.10344827586206896,0,"['books.google.com', 'books.google.com', 'douzelage.org', 'douzelage.org', 'www.rockefellerfoundation.org']",694273,Allow all users (no expiry set),44192,31 May 2004,Stan Shebs ,745,0,2004-05-31,2004-05,2004
602,602,Culture of Bangladesh,https://en.wikipedia.org/wiki/Culture_of_Bangladesh,10,0,[],[],8,0,0,2,0,0,0,0.8,0.0,0.2,0.0,0.0,0.8,0,"['www.nerdygaga.com', 'bdnews24.com', 'whc.unesco.org', 'whc.unesco.org', 'www.unesco.org', 'ich.unesco.org', 'www.unesco.org', 'whc.unesco.org', 'www.unesco.org', 'en.banglapedia.org']",1893597,Allow all users (no expiry set),32619,16 May 2005,Ragib ,1017,4,2005-05-16,2005-05,2005
603,603,Culture of Paris,https://en.wikipedia.org/wiki/Culture_of_Paris,21,1,"['10.1080/01615441003729945', None, None]",[[' historical methods']],0,0,0,6,0,0,14,0.0,0.0,0.2857142857142857,0.047619047619047616,0.0,0.047619047619047616,1,"['www.paris.location-guides.com', 'cnn.com', 'www.youtube.com', 'www.franceway.com', 'www.languagemonitor.com', 'www.youtube.com', [' historical methods']]",24194247,Allow all users (no expiry set),26226,2 September 2009,Caspian blue ,272,0,2009-09-02,2009-09,2009
604,604,Potes,https://en.wikipedia.org/wiki/Potes,1,0,[],[],0,0,0,1,0,0,0,0.0,0.0,1.0,0.0,0.0,0.0,0,['www.elpais.com'],35842677,Allow all users (no expiry set),12125,16 May 2012,Calen11 ,67,0,2012-05-16,2012-05,2012
605,605,Gaza City,https://en.wikipedia.org/wiki/Gaza_City,208,1,"['10.2307/601117', None, None]",[[' journal of the american oriental society ']],26,11,0,68,0,0,106,0.125,0.052884615384615384,0.3269230769230769,0.004807692307692308,0.0,0.18269230769230768,1,"['www.mfa.gov', 'www.pcbs.gov', 'www.pcbs.gov', 'www.pcbs.gov', 'www.pcbs.gov', 'webarchive.loc.gov', 'www.mohe.gov', 'www.pcbs.gov', 'www.pcbs.gov', 'www.pcbs.gov', 'www.gaza.gov', 'books.google.com', 'books.google.com', 'www.thisweekinpalestine.com', 'www.cbsnews.com', 'books.google.com', 'www.thisweekinpalestine.com', 'topics.nytimes.com', 'www.palestineremembered.com', 'books.google.com', 'books.google.com', 'www.com', 'www.usatoday.com', 'www.linkedin.com', 'translate.google.com', 'books.google.com', 'www.palestineremembered.com', 'nytimes.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.bbc.com', 'www.jewishencyclopedia.com', 'books.google.com', 'books.google.com', 'weather.msn.com', 'www.timeanddate.com', 'www.haaretz.com', 'books.google.com', 'books.google.com', 'www.thisweekinpalestine.com', 'www.palestineremembered.com', 'edition.cnn.com', 'books.google.com', 'books.google.com', 'books.google.com', 'extras.springer.com', 'books.google.com', 'books.google.com', 'www.thisweekinpalestine.com', 'books.google.com', 'books.google.com', 'www.jpost.com', 'uk.reuters.com', 'www.elperiodicoextremadura.com', 'www.nytimes.com', 'www.washingtonpost.com', 'www.nytimes.com', 'www.thisweekinpalestine.com', 'www.rsssf.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.csmonitor.com', 'www.palestinechronicle.com', 'books.google.com', 'www.palestineremembered.com', 'books.google.com', 'books.google.com', 'translate.google.com', 'www.google.com', 'www.worldstadia.com', 'books.google.com', 'www.jpost.com', 'books.google.com', 'translate.google.com', 'www.businessweek.com', 'www.haaretz.com', 'mediciconafrica.altervista.org', 'www.biblelands.org', 'www.mogaza.org', 'www.mogaza.org', 'www.ochaopt.org', 'www.mogaza.org', 'gisha.org', 'www.mogaza.org', 'www.english.imjnet.org', 'www.palestinecostumearchive.org', 'merip.org', 'web.nli.org', 'www.mogaza.org', 'www.mogaza.org', 'www.ochaopt.org', 'www.mogaza.org', 'www.npr.org', 'www.passia.org', 'www.christusrex.org', 'www.dci-pal.org', 'www.archnet.org', 'www.mogaza.org', 'www.cwgc.org', 'www.jewishvirtuallibrary.org', 'www.mogaza.org', 'www.globalsecurity.org', [' journal of the american oriental society ']]",55387,Require administrator access (no expiry set),115057,7 June 2002,Fredbauder ,2923,0,2002-06-07,2002-06,2002
606,606,Culture of Syria,https://en.wikipedia.org/wiki/Culture_of_Syria,22,0,[],[],1,0,0,5,0,0,16,0.045454545454545456,0.0,0.22727272727272727,0.0,0.0,0.045454545454545456,0,"['books.google.com', 'poemhunter.com', 'www.traditionalarabicmusic.com', 'www.newser.com', 'books.google.com', 'ocasia.org']",6020626,Allow all users (no expiry set),21096,18 July 2006,Kruckenberg.1 ,127,0,2006-07-18,2006-07,2006
607,607,Piacenza,https://en.wikipedia.org/wiki/Piacenza,22,0,[],[],1,1,0,3,0,0,17,0.045454545454545456,0.045454545454545456,0.13636363636363635,0.0,0.0,0.09090909090909091,0,"['ftp.atdd.noaa.gov', 'www.nytimes.com', 'www.com', 'www.piacenza-s-iano.climatemps.com', 'climaintoscana.altervista.org']",240090,Allow all users (no expiry set),38833,4 June 2003,80.180.128.130 ,781,1,2003-06-04,2003-06,2003
608,608,Ioannina,https://en.wikipedia.org/wiki/Ioannina,95,3,"['10.12681/eadd/12856', '10.1007/s11192-009-0048-4', '10.1017/s0003598x00059421', None, None, None, None, None, None]","[['didaktorika.gr', 'πανεπιστήμιο ιωαννίνων. σχολή φιλοσοφική. τμήμα ιστορίας και αρχαιολογίας. τομέας ιστορίας νεώτερων χρόνων'], ['scientometrics', 'scientometrics '], ['antiquity']]",5,1,0,33,0,0,53,0.05263157894736842,0.010526315789473684,0.3473684210526316,0.031578947368421054,0.0,0.09473684210526316,3,"['www.epirus.gov', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'travelioannina.com', 'apnews.com', 'edwardvictor.com', 'travelioannina.com', 'travelioannina.com', 'books.google.com', 'books.google.com', 'www.limassolmunicipal.com', 'www.thenationalherald.com', 'books.google.com', 'www.leidenranking.com', 'books.google.com', 'travelioannina.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'travelioannina.com', 'travelioannina.com', 'books.google.com', 'books.google.com', 'books.google.com', 'travelioannina.com', 'travelioannina.com', 'www.highbeam.com', 'www.timeshighereducation.com', 'www.travelioannina.com', 'books.google.com', 'travelioannina.com', 'www.jta.org', 'www.yadvashem.org', 'www.kkjsm.org', 'archive.adl.org', 'www.kkjsm.org', ['didaktorika.gr', 'πανεπιστήμιο ιωαννίνων. σχολή φιλοσοφική. τμήμα ιστορίας και αρχαιολογίας. τομέας ιστορίας νεώτερων χρόνων'], ['scientometrics', 'scientometrics '], ['antiquity']]",302624,Require autoconfirmed or confirmed access (no expiry set),81680,22 August 2003,195.242.150.176 ,1815,2,2003-08-22,2003-08,2003
609,609,East Frisia,https://en.wikipedia.org/wiki/East_Frisia,11,0,[],[],0,0,0,3,0,0,8,0.0,0.0,0.2727272727272727,0.0,0.0,0.0,0,"['www.britannica.com', 'www.nytimes.com', 'www.britannica.com']",146789,Allow all users (no expiry set),23175,13 November 2002,Olivier ,351,0,2002-11-13,2002-11,2002
610,610,"Crema, Lombardy","https://en.wikipedia.org/wiki/Crema,_Lombardy",4,0,[],[],0,0,0,1,0,0,3,0.0,0.0,0.25,0.0,0.0,0.0,0,['www.nytimes.com'],2252238,Allow all users (no expiry set),12727,17 July 2005,Mario Ferretti ,247,1,2005-07-17,2005-07,2005
611,611,Taranto,https://en.wikipedia.org/wiki/Taranto,46,0,[],[],3,0,0,15,0,1,27,0.06521739130434782,0.0,0.32608695652173914,0.0,0.0,0.06521739130434782,0,"['books.google.com', 'books.google.com', 'www.worldportsource.com', 'www.com', 'www.wallpaper.com', 'travelgrove.com', 'prolocoditaranto.wordpress.com', 'www.collinsdictionary.com', 'www.reuters.com', 'books.google.com', 'nobledynasty.com', 'www.imdb.com', 'ilcortiledeimelograni.wordpress.com', 'en.oxforddictionaries.com', 'italythisway.com', 'climaintoscana.altervista.org', 'phys.org', 'www.archeotaranto.altervista.org']",56148,Allow all users (no expiry set),51906,11 June 2002,Panairjdde~enwiki ,1254,4,2002-06-11,2002-06,2002
612,612,"Shaki, Azerbaijan","https://en.wikipedia.org/wiki/Shaki,_Azerbaijan",62,0,[],[],12,7,0,13,0,0,30,0.1935483870967742,0.11290322580645161,0.20967741935483872,0.0,0.0,0.3064516129032258,0,"['sheki-ih.gov', 'www.arxkom.gov', 'www.sheki-ih.gov', 'sheki-ih.gov', 'sheki-ih.gov', 'ensiklopediya.gov', 'www.mincom.gov', 'azerbaijan24.com', 'www.bostonglobe.com', 'issuu.com', 'azer.com', 'azer.com', 'gundelik-baku.com', 'varandej.livejournal.com', 'www.fallingrain.com', 'narinqala.com', 'www.orexca.com', 'books.google.com', 'guidepicker.com', 'books.google.com', 'en.unesco.org', 'lib.aliyev-heritage.org', 'whc.unesco.org', 'lib.aliyev-heritage.org', 'lib.aliyev-heritage.org', 'azadlig.org', 'iranicaonline.org', 'archnet.org', 'heydar-aliyev-foundation.org', 'www.worldcat.org', 'www.iranicaonline.org', 'www.azerembassy-kuwait.org']",1070302,Allow all users (no expiry set),38684,15 October 2004,Amiroff ,588,0,2004-10-15,2004-10,2004
613,613,Vercelli,https://en.wikipedia.org/wiki/Vercelli,6,0,[],[],1,0,0,0,0,0,5,0.16666666666666666,0.0,0.0,0.0,0.0,0.16666666666666666,0,['www.jewishitaly.org'],726056,Allow all users (no expiry set),13482,14 June 2004,Vanished user 1234567890 ,319,0,2004-06-14,2004-06,2004
614,614,Mangalorean Catholics,https://en.wikipedia.org/wiki/Mangalorean_Catholics,335,2,"['10.1007/bf00183519', '10.1515/ijsl.1978.16.77', None, None, None, None]","[[' [https'], [' international journal of the sociology of language']]",8,0,0,118,0,0,207,0.023880597014925373,0.0,0.3522388059701492,0.005970149253731343,0.0,0.029850746268656716,2,"['www.mangaloretoday.com', 'books.google.com', 'www.daijiworld.com', 'books.google.com', 'www.konkanicatholics.com', 'articles.timesofindia.indiatimes.com', 'books.google.com', 'www.daijiworld.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.konkanisongbook.com', 'books.google.com', 'books.google.com', 'hindu.com', 'hindu.com', '2fwww.daijiworld.com', 'www.hindu.com', 'books.google.com', 'books.google.com', '2fwww.daijiworld.com', 'books.google.com', 'www.geocities.com', 'www.daijiworld.com', 'books.google.com', 'www.hindu.com', 'www.hindu.com', 'books.google.com', 'www.daijiworld.com', 'books.google.com', 'www.ethnologue.com', 'www.daijiworld.com', '2fwww.mangalorean.com', 'dnaindia.com', 'books.google.com', 'mangalorean.com', 'books.google.com', 'books.google.com', 'www.khaasbaat.com', 'books.google.com', 'books.google.com', 'www.daijiworld.com', 'books.google.com', 'books.google.com', 'www.hindu.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.hindu.com', 'expressindia.indianexpress.com', 'daijiworld.com', 'books.google.com', 'books.google.com', 'www.daijiworld.com', 'books.google.com', 'books.google.com', '2fwww.daijiworld.com', 'books.google.com', 'books.google.com', '2fwww.daijiworld.com', 'books.google.com', 'www.konkanifoundation.com', '2fwww.daijiworld.com', 'www.hindu.com', 'books.google.com', 'resources.metapress.com', 'mangalorecatholicsyd.com', 'books.google.com', 'www.hinduonnet.com', 'www.daijiworld.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', '2fwww.daijiworld.com', 'www.hindu.com', 'www.daijiworld.com', 'www.daijiworld.com', 'www.indianexpress.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.daijiworld.com', 'books.google.com', 'www.daijiworld.com', 'books.google.com', 'www.daijiworld.com', 'www.daijiworld.com', 'greatest-battles.webs.com', 'www.hindu.com', 'www.daijiworld.com', 'books.google.com', 'www.daijiworld.com', 'www.daijiworld.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', '2fwww.daijiworld.com', 'www.daijiworld.com', '2fwww.mangaloretoday.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.daijiworld.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.goakonkaniakademi.org', 'www.dioceseofmangalore.org', 'stjosephseminary.org', 'quilondiocese.org', 'www.dioceseofmangalore.org', 'kcamumbai.org', 'www.mcaqatar.org', 'www.verapolyarchdiocese.org', [' [https'], [' international journal of the sociology of language']]",5474046,Allow all users (no expiry set),155712,8 June 2006,Jesuvera ,3982,3,2006-06-08,2006-06,2006
615,615,Brindisi,https://en.wikipedia.org/wiki/Brindisi,29,1,"['10.1515/9783110815931.31', None, None]",[['de gruyter mouton']],0,0,0,2,0,0,26,0.0,0.0,0.06896551724137931,0.034482758620689655,0.0,0.034482758620689655,1,"['allcorfu.com', 'wtatennis.com', ['de gruyter mouton']]",392267,Allow all users (no expiry set),52429,7 December 2003,Szopen ,610,0,2003-12-07,2003-12,2003
616,616,Żary,https://en.wikipedia.org/wiki/%C5%BBary,11,0,[],[],0,2,0,1,0,0,8,0.0,0.18181818181818182,0.09090909090909091,0.0,0.0,0.18181818181818182,0,"['stat.gov', 'www.gov', 'promienzary.com']",386902,Allow all users (no expiry set),24928,4 December 2003,Caius2ga ,213,4,2003-12-04,2003-12,2003
617,617,Erzurum,https://en.wikipedia.org/wiki/Erzurum,49,0,[],[],3,2,0,7,0,0,37,0.061224489795918366,0.04081632653061224,0.14285714285714285,0.0,0.0,0.10204081632653061,0,"['www.mgm.gov', '2009-2017.state.gov', 'books.google.com', 'books.google.com', 'erzurumguide.com', 'www.post-gazette.com', 'www.todayszaman.com', 'en.mehrnews.com', 'www.turkishpress.com', 'www.gcatholic.org', 'dergipark.org', 'archnet.org']",966195,Require autoconfirmed or confirmed access (no expiry set),41165,7 September 2004,Altenmann ,1468,4,2004-09-07,2004-09,2004
618,618,Tamil Jain,https://en.wikipedia.org/wiki/Tamil_Jain,37,0,[],[],2,0,0,15,0,0,20,0.05405405405405406,0.0,0.40540540540540543,0.0,0.0,0.05405405405405406,0,"['books.google.com', 'books.google.com', 'www.msn.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.newindianexpress.com', 'www.jainheritagecentres.com', 'akalanka-educational-trust.com', 'www.thehindu.com', 'books.google.com', 'www.thehindu.com', 'www.mustseeindia.com', 'www.jainworld.com', 'www.thenewsminute.com', 'www.tamiljains.org', 'jainsamaj.org']",665040,Allow all users (no expiry set),34543,19 May 2004,203.200.38.83 ,698,4,2004-05-19,2004-05,2004
619,619,Al-Karak,https://en.wikipedia.org/wiki/Al-Karak,49,0,[],[],2,0,0,6,0,0,41,0.04081632653061224,0.0,0.12244897959183673,0.0,0.0,0.04081632653061224,0,"['books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.ucc.org', 'babel.hathitrust.org']",307576,Allow all users (no expiry set),26476,30 August 2003,65.93.25.11 ,534,2,2003-08-30,2003-08,2003
620,620,Malatya,https://en.wikipedia.org/wiki/Malatya,46,1,[],[],6,3,0,10,0,0,26,0.13043478260869565,0.06521739130434782,0.21739130434782608,0.021739130434782608,0.0,0.21739130434782608,0,"['www.mgm.gov', 'www.malatya.gov', 'www.resmigazete.gov', 'malatyahaber.com', 'books.google.com', 'books.google.com', 'books.google.com', 'malatyaguncel.com', 'www.2theadvocate.com', 'books.google.com', 'www.milliyet.com', 'books.google.com', 'www.yenisafak.com', 'www.iranicaonline.org', 'www.jstor.org', 'www.malatyatso.org', 'en.wikisource.org', 'www.wdl.org', 'remacle.org']",1291890,Allow all users (no expiry set),41846,17 December 2004,Llywrch ,1012,2,2004-12-17,2004-12,2004
621,621,Qabala,https://en.wikipedia.org/wiki/Qabala,43,0,[],[],3,14,0,9,0,0,17,0.06976744186046512,0.32558139534883723,0.20930232558139536,0.0,0.0,0.3953488372093023,0,"['www.qebele-ih.gov', 'www.mct.gov', 'www.qebele-ih.gov', 'www.qebele-ih.gov', 'www.qebele-ih.gov', 'www.qebele-ih.gov', 'www.qebele-ih.gov', 'www.qebele-ih.gov', 'www.qebele-ih.gov', 'www.qebele-ih.gov', 'www.qebele-ih.gov', 'ftp.atdd.noaa.gov', 'www.mct.gov', 'www.mfa.gov', 'azer.com', 'qebelewelcomesyou.wordpress.com', 'www.aspiwinery.com', 'www.advantour.com', 'www.thebusinessyear.com', 'www.thebusinessyear.com', 'beltmannpianos-azerbaijan.com', 'www.booking.com', 'gilanpianos.com', 'qabala.aztelekom.org', 'www.belediyye.org', 'www.turksam.org']",2813530,Allow all users (no expiry set),24093,2 October 2005,Golbez ,316,1,2005-10-02,2005-10,2005
622,622,Hatay Province,https://en.wikipedia.org/wiki/Hatay_Province,41,0,[],[],4,6,0,20,0,0,11,0.0975609756097561,0.14634146341463414,0.4878048780487805,0.0,0.0,0.24390243902439024,0,"['kutuphane.tuik.gov', 'data.tuik.gov', 'parliament.gov', 'www.mgm.gov', 'biruni.tuik.gov', 'www.hataykulturturizm.gov', 'books.google.com', 'books.google.com', 'books.google.com', 'hurriyet.com', 'www.bbc.com', 'books.google.com', 'books.google.com', 'www.turkishpress.com', 'www.historyoftruth.com', 'books.google.com', 'books.google.com', 'www.radikal.com', 'books.google.com', 'www.jpost.com', 'books.google.com', 'www.turkishdailynews.com', 'hurarsiv.hurriyet.com', 'www.todayszaman.com', 'books.google.com', 'books.google.com', 'bianet.org', 'www.jstor.org', 'culturalsurvival.org', 'carnegieendowment.org']",403424,Allow all users (no expiry set),45869,15 December 2003,141.156.44.81 ,1113,4,2003-12-15,2003-12,2003
623,623,History of West Africa,https://en.wikipedia.org/wiki/History_of_West_Africa,256,55,"['10.1017/s0021853700000475', '10.1086/201079', '10.1080/13629387.2011.635450', '10.1023/a:1021666919678', '10.1093/hmg/ddab004', '10.1093/acrefore/9780190277734.013.137', '10.1016/j.ajhg.2019.02.007', '10.1016/j.jasrep.2020.102658', '10.2307/1166259', '10.1126/sciadv.aax5097', '10.15184/aqy.2017.30', '10.1093/acrefore/9780190854584.013.66', '10.1017/s0003598x00062840', '10.1111/j.1468-0289.2011.00627.x', '10.1016/j.nimb.2007.04.086', '10.1017/s0021853700009981', '10.1002/oa.716', '10.1093/acrefore/9780190277734.013.148', '10.1093/acrefore/9780190277734.013.285', '10.1098/rspb.2018.2288', '10.1111/ahg.12040', '10.1017/s0021853700023252', None, '10.1093/gbe/evv118', '10.1007/s10963-009-9030-6', '10.1017/s0021853700025949', '10.1080/0067270x.2012.707470', '10.4000/etudesafricaines.16965', '10.1016/j.crte.2009.04.005', '10.1016/j.ajhg.2009.05.001', '10.1386/ijia.6.1.97_1', None, '10.1098/rsos.180543', '10.1016/j.ajhg.2018.02.003', '10.1162/afar_a_00515', '10.1016/j.jas.2011.09.005', '10.1007/s12520-021-01293-5', '10.1080/21505594.2020.1809963', '10.1007/s00334-003-0016-5', '10.1038/s41598-020-79418-4', '10.1002/humu.9469', '10.2218/jls.v4i1.1682', '10.1146/annurev-genom-083117-021759', '10.1080/0067270x.2017.1393925', '10.1086/200878', '10.1002/oa.957', '10.1007/978-981-15-1614-6_10-1', '10.1534/genetics.119.302368', '10.1023/a:1015479826570', '10.3378/027.082.0402', '10.1007/s10963-019-09131-2', '10.1126/science.1172257', '10.1080/13629387.2010.486573', None, None, None, None, '33461216', None, '30827499', None, None, '32095519', None, None, None, None, None, None, None, None, None, '30963949', '25069842', None, '24089595', '26108492', None, None, None, None, None, '19500773', None, '12313941', '30225046', '29526279', None, None, '33758626', '32862777', None, '33431997', '17154278', None, '29727585', None, None, None, None, '31196864', None, '21082907', None, '19407144', None, None, None, None, None, '8117455', None, '6407493', None, None, '7015685', None, None, None, None, None, None, None, None, None, '6364581', None, None, '3786551', '4524485', None, None, None, None, None, '2694979', None, None, '6124094', '5985360', None, None, '7937602', '7549983', None, '7801626', None, None, None, None, None, None, None, '6707464', None, None, None, '2947357', None]","[['the journal of african history '], ['current anthropology'], ['the journal of north african studies '], ['african archaeological review'], ['human molecular genetics '], ['oxford university press'], ['american journal of human genetics '], ['journal of archaeological science'], ['issue', 'african studies association '], ['science advances'], ['antiquity '], ['oxford university press'], [' [[antiquity ', ' antiquity publications ltd.'], ['the economic history review '], ['nuclear instruments and methods in physics research section b'], ['the journal of african history '], ['international journal of osteoarchaeology '], ['oxford university press'], ['oxford research encyclopedias'], ['proceedings of the royal society b'], ['annals of human genetics '], ['the journal of african history '], ['sahara '], ['genome biology and evolution ', 'genome biol evol'], ['journal of world prehistory'], ['journal of african history'], ['azania'], ['cahiers d'], ['comptes rendus geoscience'], ['the american journal of human genetics'], ['international journal of islamic architecture '], [' draper fund report '], ['royal society open science ', 'royal society publishing'], ['american journal of human genetics ', 'am j hum genet.'], ['african arts'], ['journal of archaeological science '], ['archaeological and anthropological sciences '], ['virulence '], ['vegetation history and archaeobotany'], ['scientific reports '], ['human mutation'], ['journal of lithic studies'], ['annual review of genomics and human genetics '], ['azania'], ['current anthropology '], ['international journal of osteoarchaeology '], ['the handbook of mummy studies'], ['genetics '], ['[[african archaeological review'], ['human biology '], ['journal of world prehistory '], ['[[science '], ['the journal of north african studies ']]",25,8,0,60,0,0,113,0.09765625,0.03125,0.234375,0.21484375,0.0,0.34375,53,"['pdf.usaid.gov', 'aids.gov', 'www.cdc.gov', 'www.pepfar.gov', 'www.cdc.gov', 'wwwnc.cdc.gov', 'www.cdc.gov', 'www.cdc.gov', 'livescience.com', 'books.google.com', 'www.sciencedirect.com', 'search.proquest.com', 'books.google.com', 'books.google.com', 'www.newscientist.com', 'books.google.com', 'brill.com', 'www.bbc.com', 'books.google.com', 'www.cnn.com', 'findarticles.com', 'www.nytimes.com', 'www.csmonitor.com', 'search.proquest.com', 'www.bbc.com', 'translate.google.com', 'books.google.com', 'books.google.com', 'www.barakatgallery.com', 'books.google.com', 'books.google.com', 'britannica.com', 'encyclopedia.com', 'books.google.com', 'books.google.com', 'www.sciencedirect.com', 'translate.google.com', 'books.google.com', 'www.sciencedaily.com', 'translate.google.com', 'books.google.com', 'www.bbc.com', 'www.newscientist.com', 'translate.google.com', 'www.thoughtco.com', 'translate.google.com', 'books.google.com', 'africamasterweb.com', 'books.google.com', 'books.google.com', 'encyclopedia.com', 'genographic.nationalgeographic.com', 'www.hamillgallery.com', 'books.google.com', 'thinkafricapress.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.insidejustice.com', 'findarticles.com', 'books.google.com', 'oxfordre.com', 'books.google.com', 'genographic.nationalgeographic.com', 'www.dddmag.com', 'books.google.com', 'historyguy.com', 'books.google.com', 'blackpast.org', 'science.sciencemag.org', 'onafrica.org', 'unesdoc.unesco.org', 'www.publicanthropology.org', 'whc.unesco.org', '2fwhc.unesco.org', 'www.conserveafrica.org', 'advances.sciencemag.org', 'www.metmuseum.org', 'science.sciencemag.org', '2fwhc.unesco.org', '2fwhc.unesco.org', 'whc.unesco.org', 'www.ijhonline.org', 'science.sciencemag.org', '2fwhc.unesco.org', 'advances.sciencemag.org', 'whc.unesco.org', 'www.tagant.org', 'www.unaids.org', 'www.worldhistory.org', 'science.sciencemag.org', 'www.africabib.org', 'whc.unesco.org', ['the journal of african history '], ['current anthropology'], ['the journal of north african studies '], ['african archaeological review'], ['human molecular genetics '], ['oxford university press'], ['american journal of human genetics '], ['journal of archaeological science'], ['issue', 'african studies association '], ['science advances'], ['antiquity '], ['oxford university press'], [' [[antiquity ', ' antiquity publications ltd.'], ['the economic history review '], ['nuclear instruments and methods in physics research section b'], ['the journal of african history '], ['international journal of osteoarchaeology '], ['oxford university press'], ['oxford research encyclopedias'], ['proceedings of the royal society b'], ['annals of human genetics '], ['the journal of african history '], ['sahara '], ['genome biology and evolution ', 'genome biol evol'], ['journal of world prehistory'], ['journal of african history'], ['azania'], ['cahiers d'], ['comptes rendus geoscience'], ['the american journal of human genetics'], ['international journal of islamic architecture '], [' draper fund report '], ['royal society open science ', 'royal society publishing'], ['american journal of human genetics ', 'am j hum genet.'], ['african arts'], ['journal of archaeological science '], ['archaeological and anthropological sciences '], ['virulence '], ['vegetation history and archaeobotany'], ['scientific reports '], ['human mutation'], ['journal of lithic studies'], ['annual review of genomics and human genetics '], ['azania'], ['current anthropology '], ['international journal of osteoarchaeology '], ['the handbook of mummy studies'], ['genetics '], ['[[african archaeological review'], ['human biology '], ['journal of world prehistory '], ['[[science '], ['the journal of north african studies ']]",2435657,Allow all users (no expiry set),181707,12 August 2005,Dvyost ,1143,0,2005-08-12,2005-08,2005
624,624,"Ávila, Spain","https://en.wikipedia.org/wiki/%C3%81vila,_Spain",28,1,[],[],1,0,0,8,0,0,18,0.03571428571428571,0.0,0.2857142857142857,0.03571428571428571,0.0,0.07142857142857142,0,"['viajardescubriendo.com', 'www.youtube.com', 'www.avilaturismo.com', 'www.youtube.com', 'centrodeestudiosabulenses.blogia.com', 'www.collinsdictionary.com', 'books.google.com', 'periodicocorreo.com', 'www.patrimoniocastillayleon.org']",394589,Allow all users (no expiry set),33299,9 December 2003,Pfortuny ,633,2,2003-12-09,2003-12,2003
625,625,Grosseto,https://en.wikipedia.org/wiki/Grosseto,1,0,[],[],0,0,0,1,0,0,0,0.0,0.0,1.0,0.0,0.0,0.0,0,['www.com'],1054770,Allow all users (no expiry set),38667,10 October 2004,Bill Thayer ,389,0,2004-10-10,2004-10,2004
626,626,Culture of Portugal,https://en.wikipedia.org/wiki/Culture_of_Portugal,2,0,[],[],1,0,0,0,0,0,1,0.5,0.0,0.0,0.0,0.0,0.5,0,['www.wdl.org'],549666,Allow all users (no expiry set),56366,24 March 2004,PedroPVZ ,1039,0,2004-03-24,2004-03,2004
627,627,Płock,https://en.wikipedia.org/wiki/P%C5%82ock,56,2,"['10.5194/hess-11-1633-2007', '10.1127/0941-2948/2006/0130', None, None, None, None]","[['hydrol. earth syst. sci. '], ['meteorologische zeitschrift']]",4,4,0,3,0,0,43,0.07142857142857142,0.07142857142857142,0.05357142857142857,0.03571428571428571,0.0,0.17857142857142858,2,"['bdl.stat.gov', 'www.gov', 'bdl.stat.gov', 'www.gov', 'mostwplocku.blogspot.com', 'samgrubersjewishartmonuments.blogspot.com', 'www.eilatgordinlevitan.com', 'malachowianka.plock.org', 'www.sztetl.org', 'www.sztetl.org', 'www.sztetl.org', ['hydrol. earth syst. sci. '], ['meteorologische zeitschrift']]",74609,Allow all users (no expiry set),46493,22 August 2002,217.99.105.223 ,617,1,2002-08-22,2002-08,2002
628,628,Patras,https://en.wikipedia.org/wiki/Patras,83,0,[],[],4,3,0,9,0,1,66,0.04819277108433735,0.03614457831325301,0.10843373493975904,0.0,0.0,0.08433734939759036,0,"['dikitiellada.gov', 'dikitiellada.gov', 'ditikiellada.gov', 'translate.yandex.com', 'ditikiellda-region.com', 'ktizon.blogspot.com', 'greekreporter.com', 'intracom-telecom.com', 'www.ditikiellada-region.com', 'acciona-energia.com', 'www.ditikiellada-region.com', 'www.limassolmunicipal.com', 'www.sister-cities.org', 'www.psp.org', 'corallia.org', 'europe.anglican.org']",470691,Allow all users (no expiry set),95076,15 February 2004,Ikariotis ,2667,0,2004-02-15,2004-02,2004
629,629,Treviso,https://en.wikipedia.org/wiki/Treviso,30,0,[],[],0,1,0,8,0,0,21,0.0,0.03333333333333333,0.26666666666666666,0.0,0.0,0.03333333333333333,0,"['www.cmc.pr.gov', 'www.weatherbase.com', 'books.google.com', 'www.marcadoc.com', 'weatherbase.com', 'goodtimefortrip.com', 'www.com', 'www.com', 'www.nytimes.com']",925340,Allow all users (no expiry set),35186,24 August 2004,Waltpohl ,535,3,2004-08-24,2004-08,2004
630,630,Outline of Andhra Pradesh,https://en.wikipedia.org/wiki/Outline_of_Andhra_Pradesh,1,0,[],[],1,0,0,0,0,0,0,1.0,0.0,0.0,0.0,0.0,1.0,0,['svzoo.org'],44143246,Allow all users (no expiry set),17346,18 October 2014,AhamSarvatra ,131,0,2014-10-18,2014-10,2014
631,631,Oron people,https://en.wikipedia.org/wiki/Oron_people,50,1,"['10.2307/1156343', None, None]",[['africa']],5,1,0,22,0,0,21,0.1,0.02,0.44,0.02,0.0,0.14,1,"['www.nipost.gov', 'books.google.com', 'www.abebooks.com', 'www.premiumtimesng.com', 'books.google.com', 'www.manpower.com', 'akwaibomcelebrates.com', 'books.google.com', 'www.premiumtimesng.com', 'books.google.com', 'the-nigeria.com', 'www.artkhade.com', 'www.abebooks.com', 'nm.onlinenigeria.com', 'www.abebooks.com', 'books.google.com', 'books.google.com', 'www.city-facts.com', 'www.abebooks.com', 'dailyindependentnig.com', 'nationalnewstrack.com', 'www.abebooks.com', 'www.abebooks.com', 'www.nassnig.org', 'www.nassnig.org', 'www.waado.org', 'www.ambazoniagov.org', 'www.jstor.org', ['africa']]",20784669,Allow all users (no expiry set),88110,20 December 2008,Utibe10 ,510,5,2008-12-20,2008-12,2008
632,632,Maniots,https://en.wikipedia.org/wiki/Maniots,112,1,"['10.1038/ejhg.2017.18', '28272534', '5437898']",[['european journal of human genetics']],3,0,0,2,0,0,106,0.026785714285714284,0.0,0.017857142857142856,0.008928571428571428,0.0,0.03571428571428571,1,"['books.google.com', 'books.google.com', 'www.mani.org', 'mani.org', 'www.mani.org', ['european journal of human genetics']]",2266821,Allow all users (no expiry set),89822,19 July 2005,64.136.27.225 ,1403,1,2005-07-19,2005-07,2005
633,633,Jammu division,https://en.wikipedia.org/wiki/Jammu_division,114,0,[],[],1,24,0,71,0,0,18,0.008771929824561403,0.21052631578947367,0.6228070175438597,0.0,0.0,0.21929824561403508,0,"['www.censusindia.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'censusindia.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'censusindia.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'censusindia.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'censusindia.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'censusindia.gov', 'www.censusindia.gov', 'www.censusindia.gov', 'censusindia.gov', 'books.google.com', 'www.dailyexcelsior.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.dailyexcelsior.com', 'books.google.com', 'www.dailyexcelsior.com', 'books.google.com', 'www.dailyexcelsior.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.dailyexcelsior.com', 'www.dailyexcelsior.com', 'www.bhaderwah.com', 'www.indictoday.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thehindu.com', 'books.google.com', 'www.dailyexcelsior.com', 'www.outlookindia.com', 'www.firstpost.com', 'books.google.com', 'books.google.com', 'books.google.com', 'economictimes.indiatimes.com', 'books.google.com', 'www.news18.com', 'books.google.com', 'www.jammu-kashmir.com', 'www.dailyexcelsior.com', 'books.google.com', 'risingkashmir.com', 'www.tribuneindia.com', 'books.google.com', 'books.google.com', 'www.dailyexcelsior.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.dailyexcelsior.com', 'www.dailyexcelsior.com', 'www.dailyexcelsior.com', 'books.google.com', 'books.google.com', 'www.tribuneindia.com', 'www.livemint.com', 'books.google.com', 'books.google.com', 'www.dailyexcelsior.com', 'outlookindia.com', 'books.google.com', 'books.google.com', 'economictimes.indiatimes.com', 'books.google.com', 'books.google.com', 'www.dailyexcelsior.com', 'books.google.com', 'books.google.com', 'www.orfonline.org']",43066131,Allow all users (no expiry set),97262,16 March 2004,202.138.119.193 ,1530,4,2004-03-16,2004-03,2004
634,634,Metsovo,https://en.wikipedia.org/wiki/Metsovo,14,0,[],[],0,0,0,4,0,0,10,0.0,0.0,0.2857142857142857,0.0,0.0,0.0,0,"['books.google.com', 'books.google.com', 'books.google.com', 'books.google.com']",756618,Allow all users (no expiry set),36156,26 June 2004,24.184.180.73 ,349,0,2004-06-26,2004-06,2004
635,635,Volos,https://en.wikipedia.org/wiki/Volos,32,3,"['10.1080/20548923.2018.1427182', '10.1093/acref/9780199545568.001.0001', None, None, None, None]","[[' star', (' kastro palaia settlement', ' settlement', 'settlement', 'v')], [' oxford university press ']]",0,0,0,3,0,0,26,0.0,0.0,0.09375,0.09375,0.0,0.09375,2,"['macedonia.kroraina.com', 'books.google.com', 'books.google.com', [' star', (' kastro palaia settlement', ' settlement', 'settlement', 'v')], [' oxford university press ']]",422886,Allow all users (no expiry set),40484,6 January 2004,Sofos ,1555,3,2004-01-06,2004-01,2004
636,636,Maldivians,https://en.wikipedia.org/wiki/Maldivians,35,1,"['10.1002/ajpa.22256', '23526367', '3652038']",[['[[american journal of physical anthropology']],0,5,0,22,0,0,7,0.0,0.14285714285714285,0.6285714285714286,0.02857142857142857,0.0,0.17142857142857143,1,"['statisticsmaldives.gov', 'www.dfat.gov', 'presidencymaldives.gov', 'statisticsmaldives.gov', 'artgallery.gov', 'www.dhivehiobserver.com', 'webcache.googleusercontent.com', 'sinhalaya.com', 'minivannewsarchive.com', 'www.ethnologue.com', 'afp.google.com', 'books.google.com', 'maldivesmission.com', 'books.google.com', 'www.maldives-ethnography.com', 'www.islamkalender.com', 'everyculture.com', 'haveeru.com', 'policyresearchgroup.com', 'maldivesroyalfamily.com', 'cache:kekph3it1ssj:lt-lt.facebook.com', 'books.google.com', 'www.mathaaran.com', 'books.google.com', 'maldives-ancestry.blogspot.com', 'www.maldivesculture.com', 'www.maldivesroyalfamily.com', ['[[american journal of physical anthropology']]",23582208,Allow all users (no expiry set),55738,12 July 2009,Deviathan~enwiki ,582,1,2009-07-12,2009-07,2009
637,637,The Fisherman's Cot,https://en.wikipedia.org/wiki/The_Fisherman%27s_Cot,8,0,[],[],0,0,0,3,0,0,5,0.0,0.0,0.375,0.0,0.0,0.0,0,"['books.google.com', 'books.google.com', 'books.google.com']",30050820,Allow all users (no expiry set),5167,14 December 2010,Dr. Blofeld ,53,1,2010-12-14,2010-12,2010
638,638,Culture of Mangalorean Catholics,https://en.wikipedia.org/wiki/Culture_of_Mangalorean_Catholics,106,0,[],[],1,0,0,55,0,0,50,0.009433962264150943,0.0,0.5188679245283019,0.0,0.0,0.009433962264150943,0,"['books.google.com', 'books.google.com', 'www.hinduonnet.com', 'www.hinduonnet.com', 'greatest-battles.webs.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.hindu.com', 'www.daijiworld.com', 'www.hindu.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.hinduonnet.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.daijiworld.com', 'books.google.com', 'books.google.com', 'www.konkanifoundation.com', 'books.google.com', 'books.google.com', 'www.daijiworld.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'richardcrasta.com', 'books.google.com', 'books.google.com', 'www.hinduonnet.com', 'books.google.com', 'books.google.com', 'books.google.com', 'daijiworld.com', 'books.google.com', 'www.hinduonnet.com', 'www.daijiworld.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.daijiworld.com', 'books.google.com', 'books.google.com', 'www.ethnologue.com', 'www.theindiancatholic.com', 'www.konkanifoundation.com', 'www.goakonkaniakademi.org']",19087356,Allow all users (no expiry set),46930,29 August 2008,Kensplanet ,126,0,2008-08-29,2008-08,2008
639,639,Palencia,https://en.wikipedia.org/wiki/Palencia,10,0,[],[],0,0,0,0,0,0,10,0.0,0.0,0.0,0.0,0.0,0.0,0,[],616252,Allow all users (no expiry set),26827,24 April 2004,Montrealais ,414,0,2004-04-24,2004-04,2004
640,640,Culture in Berlin,https://en.wikipedia.org/wiki/Culture_in_Berlin,65,0,[],[],8,0,0,22,0,2,35,0.12307692307692308,0.0,0.3384615384615385,0.0,0.0,0.12307692307692308,0,"['www.observer.com', 'www.metrotimes.com', 'www.businessweek.com', 'germancorner.com', 'www.scc-events.com', 'www.newcolonist.com', 'travel.nytimes.com', 'gaytravel.about.com', 'www.washingtonpost.com', 'expatica.com', 'www.lollapaloozade.com', 'travel2.nytimes.com', 'www.slowtravelberlin.com', 'www.fifa.com', 'www.fifa.com', 'www.expatica.com', 'www.culturekiosque.com', 'www.passportmagazine.com', 'www.nytimes.com', 'blogs.bettor.com', 'www.theage.com', 'www.observer.com', 'www.metropolis2005.org', 'www.metropolis2005.org', 'thomaspainescorner.org', 'whc.unesco.org', 'www.olympic.org', 'www.berlin2009.org', 'www.europeanfilmacademy.org', 'www.germanfoods.org']",34638621,Allow all users (no expiry set),44429,7 February 2012,FinnishDriver ,120,0,2012-02-07,2012-02,2012
641,641,Ferrara,https://en.wikipedia.org/wiki/Ferrara,69,0,[],[],4,1,0,16,0,0,48,0.057971014492753624,0.014492753623188406,0.2318840579710145,0.0,0.0,0.07246376811594203,0,"['www1.interno.gov', 'www.britannica.com', 'servizi.com', 'www.ferrarainfo.com', 'books.google.com', 'www.com', 'books.google.com', 'www.nytimes.com', 'emiliaromagnaturismo.com', 'books.google.com', 'www.thestadiumbusiness.com', 'books.google.com', 'www.ft.com', 'www.com', 'emiliaromagnaturismo.com', 'www.tabletmag.com', 'www.com', 'www.napoleon-series.org', 'www.napoleon-series.org', 'www.napoleon-series.org', 'www.napoleon-series.org']",45846,Allow all users (no expiry set),52353,24 March 2002,Gianfranco ,916,0,2002-03-24,2002-03,2002
642,642,Chandannagar,https://en.wikipedia.org/wiki/Chandannagar,26,0,[],[],3,4,0,14,0,0,5,0.11538461538461539,0.15384615384615385,0.5384615384615384,0.0,0.0,0.2692307692307692,0,"['censusindia.gov', 'mea.gov', 'policewb.gov', 'www.wbpspm.gov', 'www.wbtrafficpolice.com', 'www.telegraphindia.com', 'timesofindia.indiatimes.com', 'www.thehindu.com', 'www.telegraphindia.com', 'www.telegraphindia.com', 'heritagechandernagoreblog.wordpress.com', 'timesofindia.indiatimes.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.livemint.com', 'rangandatta.wordpress.com', 'books.google.com', 'www.thehindu.com', 'en.banglapedia.org', 'www.gutenberg.org', 'www.gutenberg.org']",1470431,Allow all users (no expiry set),46205,5 February 2005,Tom Radulovich ,1092,1,2005-02-05,2005-02,2005
643,643,Parma,https://en.wikipedia.org/wiki/Parma,16,0,[],[],1,0,0,5,0,0,10,0.0625,0.0,0.3125,0.0,0.0,0.0625,0,"['www.com', 'books.google.com', 'pitoresco.com', 'www.monasterosangiovanni.com', 'books.google.com', 'www.briarpress.org']",24231,Allow all users (no expiry set),38762,30 September 2001,Trimalchio ,949,7,2001-09-30,2001-09,2001
644,644,Culture of Gujarat,https://en.wikipedia.org/wiki/Culture_of_Gujarat,22,0,[],[],0,0,0,9,0,0,13,0.0,0.0,0.4090909090909091,0.0,0.0,0.0,0,"['madhursangam.com', 'www.screenindia.com', 'www.screenindia.com', 'www.dnaindia.com', 'www.hinduismtoday.com', 'timesofindia.indiatimes.com', 'books.google.com', 'www.financialexpress.com', 'www.business-standard.com']",16568193,Allow all users (no expiry set),41678,25 March 2008,Ilikeeatingwaffles ,324,0,2008-03-25,2008-03,2008
645,645,Culture of Mongolia,https://en.wikipedia.org/wiki/Culture_of_Mongolia,24,0,[],[],7,0,0,7,0,0,10,0.2916666666666667,0.0,0.2916666666666667,0.0,0.0,0.2916666666666667,0,"['www.nytimes.com', 'www.infomongolia.com', 'money.cnn.com', 'books.google.com', 'members.aol.com', 'asianart.com', 'www.cnn.com', 'www.unesco.org', 'unesco.org', 'www.unesco.org', 'www.unesco.org', 'unesco.org', 'www.unesco.org', 'www.unesco.org']",495256,Allow all users (no expiry set),28258,29 February 2004,24.160.94.214 ,760,0,2004-02-29,2004-02,2004
646,646,Outline of Telangana,https://en.wikipedia.org/wiki/Outline_of_Telangana,4,0,[],[],0,0,0,2,0,0,2,0.0,0.0,0.5,0.0,0.0,0.0,0,"['books.google.com', 'www.newindianexpress.com']",47344138,Allow all users (no expiry set),11161,26 July 2015,Trmwikifa ,68,0,2015-07-26,2015-07,2015
647,647,List of Egyptian inventions and discoveries,https://en.wikipedia.org/wiki/List_of_Egyptian_inventions_and_discoveries,308,29,"[None, '10.1002/cncr.25553', '10.1039/b606268g', '10.2307/2973180', None, '10.1093/jss/26.2.229', '10.1016/j.nephro.2009.06.001', '10.11141/ia.42.6.3', '10.1007/s11157-007-9120-9', '10.1016/0301-0104(96)00067-5', '10.1126/science.287.5453.631', '10.2307/j.ctt21c4td4.10', '10.1080/05775132.1993.11471653', '10.2307/3209606', '10.1016/j.jvs.2014.04.056', '10.1038/s41598-021-90759-6', '10.1371/journal.pone.0144140', '10.1021/jp001460h', '10.1177/014107689608900813', '10.1007/bf02986998', '10.1016/j.jcrs.2008.11.052', '10.1016/j.jcws.2012.04.002', '10.1088/0004-637x/773/1/1', '10.1017/s0025727300028386', '10.1021/cr020689l', '10.1017/s0959774308000395', '10.2308/0148-4184.29.1.195', '10.11141/ia.42.6.5', '10.1093/oxfordhb/9780199935390.013.48', '5322341', '20960499', '17173142', None, None, None, '19617021', None, None, None, '10649992', None, None, None, '24970660', '34050218', '26679699', None, '8795503', None, '19251160', '24525756', None, '13960613', '15080722', None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, None, '8163881', '4683080', None, '1295891', None, None, '3601883', None, '1034829', None, None, None, None, None]","[['surgery '], ['cancer '], ['chemical society reviews '], [' [[the american mathematical monthly'], ['journal of archaeological science '], ['[[journal of semitic studies'], ['nephrologie '], ['internet archaeology '], ['reviews in environmental science and bio'], ['chemical physics'], ['science'], ['university college london press '], ['challenge'], [' the biblical archaeologist'], ['journal of vascular surgery'], ['scientific reports '], [' plos one'], ['the journal of physical chemistry a'], ['journal of the royal society of medicine '], ['the mathematical intelligencer '], ['journal of cataract '], [' the journal of the american college of certified wound specialists'], [' the astrophysical journal'], ['medical history'], ['chemical reviews'], [' cambridge archaeological journal'], ['accounting historians journal'], ['internet archaeology '], ['oxford handbooks online ', 'oxford university press ']]",22,1,0,93,0,0,162,0.07142857142857142,0.003246753246753247,0.30194805194805197,0.09415584415584416,0.0,0.16883116883116883,29,"['www.sis.gov', 'www.houstonspediatricdentist.com', 'www.davidensemble.com', 'www.zmescience.com', 'www.britannica.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.washingtonpost.com', 'www.historyofglass.com', 'www.tobaccopipes.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.newscientist.com', 'www.guinnessworldrecords.com', 'study.com', 'www.thrillist.com', 'www.latimes.com', 'www.themarysue.com', 'study.com', 'books.google.com', 'www.infoplease.com', 'www.newscientist.com', 'beta.theglobeandmail.com', 'egyptianmath.blogspot.com', 'eltident.com', 'worldcomp-proceedings.com', 'science.howstuffworks.com', 'books.google.com', 'helpwithbowling.com', 'www.livescience.com', 'www.si.com', 'www.msc-conf.com', 'egyptianstreets.com', 'books.google.com', 'science.howstuffworks.com', 'www.gol27.com', 'hellenicnews.com', 'time.com', 'www.history.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.pipe-maker.com', 'www.nbcnews.com', 'interestingengineering.com', 'books.google.com', 'www.boyercandies.com', 'science.howstuffworks.com', 'books.google.com', 'www.brighthubengineering.com', 'books.google.com', 'www.mrcophth.com', 'discoveringegypt.com', 'www.nytimes.com', 'scienceworld.wolfram.com', 'books.google.com', 'books.google.com', 'egyptianmath.blogspot.com', 'www.britannica.com', 'www.popularmechanics.com', 'egyptindependent.com', 'books.google.com', 'www.nytimes.com', 'www.campfiremarshmallows.com', 'books.google.com', 'www.smithsonianmag.com', 'www.upi.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.thoughtco.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'books.google.com', 'www.moundtop.com', 'books.google.com', 'books.google.com', 'www.britannica.com', 'books.google.com', 'www.upi.com', 'www.davidensemble.com', 'www.world-mysteries.com', 'egyptindependent.com', 'www.compoundchem.com', 'books.google.com', 'catchnews.com', 'delanceyplace.com', 'www.nbcnews.com', 'www.bbc.com', 'www.archaeology.org', 'www.egyptianolympic.org', 'nobelprize.org', 'www.britishmuseum.org', 'lead.org', 'www.invent.org', 'mnhs.org', 'pbs.org', 'www.asce.org', 'www.isradiology.org', 'www.npr.org', 'www.wonderopolis.org', 'www.reshafim.org', 'www.americangemsociety.org', 'www.eternalegypt.org', 'www.egyptorigins.org', 'st-takla.org', 'archaeology.org', 'english.ahram.org', 'www.cut-the-knot.org', 'www.sciencehistory.org', 'www.reshafim.org', ['surgery '], ['cancer '], ['chemical society reviews '], [' [[the american mathematical monthly'], ['journal of archaeological science '], ['[[journal of semitic studies'], ['nephrologie '], ['internet archaeology '], ['reviews in environmental science and bio'], ['chemical physics'], ['science'], ['university college london press '], ['challenge'], [' the biblical archaeologist'], ['journal of vascular surgery'], ['scientific reports '], [' plos one'], ['the journal of physical chemistry a'], ['journal of the royal society of medicine '], ['the mathematical intelligencer '], ['journal of cataract '], [' the journal of the american college of certified wound specialists'], [' the astrophysical journal'], ['medical history'], ['chemical reviews'], [' cambridge archaeological journal'], ['accounting historians journal'], ['internet archaeology '], ['oxford handbooks online ', 'oxford university press ']]",64283032,Allow all users (no expiry set),152645,15 June 2020,Mark Wagdy El-Magrisy ,433,1,2020-06-15,2020-06,2020
648,648,Vaqueiros de alzada,https://en.wikipedia.org/wiki/Vaqueiros_de_alzada,72,0,[],[],2,1,0,6,0,0,63,0.027777777777777776,0.013888888888888888,0.08333333333333333,0.0,0.0,0.041666666666666664,0,"['pubmed.ncbi.nlm.nih.gov', 'www.cervantesvirtual.com', 'issuu.com', 'www.cervantesvirtual.com', 'issuu.com', 'www.vaquerosalzadatorrestio.com', 'www.cervantesvirtual.com', 'www.semanticscholar.org', 'www.amisalas.org']",1369435,Allow all users (no expiry set),28299,7 January 2005,OldakQuill ,81,2,2005-01-07,2005-01,2005
649,649,Culture of Milan,https://en.wikipedia.org/wiki/Culture_of_Milan,33,0,[],[],5,0,0,16,0,0,12,0.15151515151515152,0.0,0.48484848484848486,0.0,0.0,0.15151515151515152,0,"['britannica.com', 'www.britannica.com', 'pasticceriacova.com', 'milan.world-guides.com', 'aboutmilan.com', 'livescience.com', 'frieze.com', 'www.americanchronicle.com', 'www.wiley.com', 'europe-cities.com', 'www.lifeinitaly.com', 'www.whatsonwhen.com', 'milan.wantedineurope.com', 'lankaramaya.com', 'languagemonitor.com', 'www.britannica.com', 'iop.org', 'orthodoxeurope.org', 'www.unipiams.org', 'newadvent.org', 'www.unipiams.org']",25477003,Allow all users (no expiry set),47897,18 December 2009,Theologiae ,219,0,2009-12-18,2009-12,2009
650,650,Culture of Hungary,https://en.wikipedia.org/wiki/Culture_of_Hungary,20,0,[],[],3,0,0,9,0,0,8,0.15,0.0,0.45,0.0,0.0,0.15,0,"['www.bbc.com', 'encyclopedia.com', 'sports-reference.com', 'herend.com', 'imdb.com', 'www.imdb.com', 'imdb.com', 'www.imdb.com', 'www.lonelyplanet.com', 'olympedia.org', 'fina.org', 'olympic.org']",869096,Allow all users (no expiry set),45839,31 July 2004,RetiredUser2 ,1347,0,2004-07-31,2004-07,2004
651,651,Culture of Pakistan,https://en.wikipedia.org/wiki/Culture_of_Pakistan,14,0,[],[],6,0,0,6,0,0,2,0.42857142857142855,0.0,0.42857142857142855,0.0,0.0,0.42857142857142855,0,"['dawn.com', 'books.google.com', 'pakistaniat.com', 'books.google.com', 'www.warc.com', 'www.dawn.com', 'www.metmuseum.org', 'whc.unesco.org', 'fao.org', 'www.theismaili.org', 'history-world.org', 'www.worldhockey.org']",1622957,Allow all users (no expiry set),31578,19 March 2005,193.220.82.125 ,2128,4,2005-03-19,2005-03,2005
652,652,Western Norway,https://en.wikipedia.org/wiki/Western_Norway,57,4,"['10.1016/0169-555x(94)90029-9', '10.1080/04353676.1967.11879749', '10.1016/s0921-8181(00)00009-6', '10.1016/0169-555x(92)90022-g', None, None, None, None, None, None, None, None]","[['[[geomorphology '], ['[[geografiska annaler'], ['[[global and planetary change'], [' [[geomorphology ']]",1,2,0,2,0,0,48,0.017543859649122806,0.03508771929824561,0.03508771929824561,0.07017543859649122,0.0,0.12280701754385964,4,"['www.cia.gov', 'state.gov', 'www.hurtigruten.com', 'ft.com', 'nobelprize.org', ['[[geomorphology '], ['[[geografiska annaler'], ['[[global and planetary change'], [' [[geomorphology ']]",1436846,Allow all users (no expiry set),77308,27 January 2005,Egil ,529,0,2005-01-27,2005-01,2005
653,653,Slobbovia,https://en.wikipedia.org/wiki/Slobbovia,0,0,[],[],0,0,0,0,0,0,0,,,,,,,0,[],3220719,Allow all users (no expiry set),55301,22 November 2005,GABaker ,270,0,2005-11-22,2005-11,2005
654,654,"Outline of Punjab, India","https://en.wikipedia.org/wiki/Outline_of_Punjab,_India",1,0,[],[],0,0,0,0,0,0,1,0.0,0.0,0.0,0.0,0.0,0.0,0,[],51466350,Allow all users (no expiry set),13212,30 August 2016,The Transhumanist ,108,0,2016-08-30,2016-08,2016
655,655,Frutigen,https://en.wikipedia.org/wiki/Frutigen,23,0,[],[],0,0,0,1,0,0,22,0.0,0.0,0.043478260869565216,0.0,0.0,0.0,0,['world.com'],4541009,Allow all users (no expiry set),25923,28 March 2006,BillC ,98,0,2006-03-28,2006-03,2006
656,656,List of Indonesian inventions and discoveries,https://en.wikipedia.org/wiki/List_of_Indonesian_inventions_and_discoveries,87,3,"['10.2307/1124435', '10.1016/s0740-0020(86)80035-1', '10.1525/aa.1987.89.2.02a00030', None, None, None, None, None, None]","[[' asian theatre journal '], ['food microbiology '], ['american anthropologist']]",5,0,0,44,0,0,35,0.05747126436781609,0.0,0.5057471264367817,0.034482758620689655,0.0,0.09195402298850575,3,"['books.google.com', 'books.google.com', 'books.google.com', 'www.1843magazine.com', 'books.google.com', 'www.theindependent.com', 'books.google.com', 'www.thejakartapost.com', 'id.berita.yahoo.com', 'www.thejakartapost.com', 'indo.com', 'books.google.com', 'www.britannica.com', 'www.kastenmarine.com', 'query.nytimes.com', 'www.bali.com', 'www.blackbeltmag.com', 'books.google.com', 'inet.detik.com', 'www.airframer.com', 'sulawesistudies.blogspot.com', 'www.beritasatu.com', 'books.google.com', 'www.ilmutekniksipil.com', 'finance.detik.com', 'www.constructionasiaonline.com', 'www.thejakartaglobe.com', 'www.thejakartapost.com', 'www.angkasa-online.com', 'papanidea.com', 'sumedangonline.com', 'www.thejakartapost.com', 'www.patentsencyclopedia.com', 'www.thejakartapost.com', 'www.thejakartapost.com', 'www.britannica.com', 'www.britannica.com', 'enviplast.com', 'www.farsidemusic.com', 'www.keganpaul.com', 'www.farsidemusic.com', 'voices.nationalgeographic.com', 'www.thejakartapost.com', 'www.thejakartapost.com', 'www.bwtp.org', 'blogs.unicef.org', 'www.insideindonesia.org', 'metmuseum.org', 'metmuseum.org', [' asian theatre journal '], ['food microbiology '], ['american anthropologist']]",43579256,Allow all users (no expiry set),60843,16 August 2014,Si Gam ,330,1,2014-08-16,2014-08,2014
657,657,Ramgarh district,https://en.wikipedia.org/wiki/Ramgarh_district,85,0,[],[],10,12,0,40,0,0,24,0.11764705882352941,0.1411764705882353,0.47058823529411764,0.0,0.0,0.25882352941176473,0,"['fossil.energy.gov', 'www.jharkhand.gov', 'www.cia.gov', '2010.census.gov', 'www.ser.indianrailways.gov', 'www.censusindia.gov', 'ccl.gov', 'www.jharkhand.gov', 'fossil.energy.gov', 'www.jharkhand.gov', 'ccl.gov', 'www.censusindia.gov', 'www.winentrance.com', 'www.jagran.com', 'www.facebook.com', 'b.com', 'www.youtube.com', 'articles.timesofindia.indiatimes.com', 'epaper.jagran.com', 'epaper.jagran.com', 'jharkhandforest.com', 'www.tatasteel.com', 'www.jagran.com', 'indianmovements.blogspot.com', 'www.jagran.com', 'www.indiamapssite.com', 'epaper.bhaskar.com', 'www.telegraphindia.com', 'www.winentrance.com', 'www.telegraphindia.com', 'indiarailinfo.com', 'www.youtube.com', 'im23-c75.kxcdn.com', 'astrobix.com', 'epaper.jagran.com', 'www.onlytravelguide.com', 'www.jagran.com', 'lawyerrlalwani.com', 'www.telegraphindia.com', 'therungtagroup.com', 'www.telegraphindia.com', 'intachranchi.com', 'www.jagran.com', 'www.livehindustan.com', 'books.google.com', 'books.google.com', 'www.jagran.com', 'epaper.jagran.com', 'im23-c75.kxcdn.com', 'www.jharkhandforest.com', 'apsramgarhcantt.com', 'im22-c75.kxcdn.com', 'www.serranchi.org', 'www.ramgarhcollege.org', 'aicc.org', 'gandhiserve.org', 'www.museumlife.org', 'www.gandhimedia.org', 'www.mkgandhi-sarvodaya.org', 'www.asiapacificpartnership.org', 'rotaryramgarh.org', 'www.mkgandhi-sarvodaya.org']",21449113,Allow all users (no expiry set),67875,8 February 2009,Ranjitsharma ,854,1,2009-02-08,2009-02,2009
658,658,Lower Assam,https://en.wikipedia.org/wiki/Lower_Assam,31,0,[],[],0,0,0,1,0,0,30,0.0,0.0,0.03225806451612903,0.0,0.0,0.0,0,['books.google.com'],25111333,Allow all users (no expiry set),24517,17 November 2009,Bhaskarbhagawati ,320,0,2009-11-17,2009-11,2009
659,659,Hunting in Romania,https://en.wikipedia.org/wiki/Hunting_in_Romania,3,0,[],[],0,0,0,0,0,0,3,0.0,0.0,0.0,0.0,0.0,0.0,0,[],20828299,Allow all users (no expiry set),29510,24 December 2008,LeonisRugitur ,428,0,2008-12-24,2008-12,2008
660,660,Umaidpur,https://en.wikipedia.org/wiki/Umaidpur,25,0,[],[],0,4,0,13,0,0,8,0.0,0.16,0.52,0.0,0.0,0.16,0,"['panchayatdirectory.gov', 'censusindia.gov', 'panchayatdirectory.gov', 'censusindia.gov', 'accuweather.com', 'indiamapped.com', 'www.bhojpuria.com', 'www.geolysis.com', 'biharandjharkhand.com', 'mapsofindia.com', 'google.com', 'geolysis.com', 'bawarchi.com', 'maps.google.com', 'distancesfrom.com', 'books.google.com', 'weather.yahoo.com']",42192517,Allow all users (no expiry set),31046,13 March 2014,Susie9 ,552,0,2014-03-13,2014-03,2014
661,661,Outline of Africa,https://en.wikipedia.org/wiki/Outline_of_Africa,0,0,[],[],0,0,0,0,0,0,0,,,,,,,0,[],16584849,Allow all users (no expiry set),18267,26 March 2008,The Transhumanist ,302,0,2008-03-26,2008-03,2008
662,662,Montagnana,https://en.wikipedia.org/wiki/Montagnana,2,0,[],[],0,0,0,0,0,0,2,0.0,0.0,0.0,0.0,0.0,0.0,0,[],1146074,Allow all users (no expiry set),10043,8 November 2004,Pumpie ,123,1,2004-11-08,2004-11,2004
663,663,Alcamo,https://en.wikipedia.org/wiki/Alcamo,151,0,[],[],3,0,0,29,0,0,119,0.019867549668874173,0.0,0.19205298013245034,0.0,0.0,0.019867549668874173,0,"['www.com', 'books.google.com', 'www.alpauno.com', 'www.com', 'www.com', 'www.com', 'www.com', 'www.com', 'www.com', 'www.com', 'books.google.com', 'www.forgottenbooks.com', 'www.com', 'www.com', 'books.google.com', 'www.com', 'www.youtube.com', 'www.com', 'www.com', 'www.com', 'www.com', 'www.com', 'www.com', 'www.com', 'www.com', 'www.gingerandtomato.com', 'www.ioamolasicilia.com', 'www.youtube.com', 'www.termelibere.com', 'arcobaleno1.altervista.org', 'climate-data.org', 'climate-data.org']",44767,Allow all users (no expiry set),99917,18 March 2002,Ik1tzo~enwiki ,1070,0,2002-03-18,2002-03,2002
664,664,Tetovo,https://en.wikipedia.org/wiki/Tetovo,45,0,[],[],2,4,0,25,0,1,13,0.044444444444444446,0.08888888888888889,0.5555555555555556,0.0,0.0,0.13333333333333333,0,"['www.stat.gov', 'tetova.gov', 'makstat.stat.gov', 'www.stat.gov', 'books.google.com', 'tetovobienale.webs.com', 'www.oup.com', 'books.google.com', 'books.google.com', 'skopje.cafebabel.com', 'books.google.com', 'www.balkantravellers.com', 'www.newsobserver.com', 'books.google.com', 'www.nytimes.com', 'books.google.com', 'www.amazon.com', 'books.google.com', 'tetova1.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.utrinski.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.balwois.com', 'www.tetovo.g3z.com', 'www.tdvia.org', 'www.ifrc.org']",1053601,Allow all users (no expiry set),53862,10 October 2004,Etz Haim ,1496,5,2004-10-10,2004-10,2004
665,665,Cuttack,https://en.wikipedia.org/wiki/Cuttack,61,1,"['10.1109/i2ct.2017.8226150', None, None]",[['2017 2nd international conference for convergence in technology ']],7,12,0,18,0,1,22,0.11475409836065574,0.19672131147540983,0.29508196721311475,0.01639344262295082,0.0,0.32786885245901637,1,"['censusindia.gov', 'www.cmccuttack.gov', 'imdpune.gov', 'paradipport.gov', 'www.rajbhavanodisha.gov', 'www.cmccuttack.gov', 'orissa.gov', 'www.cmccuttack.gov', 'imdpune.gov', 'orissa.gov', 'www.cmccuttack.gov', 'allindiaradio.gov', 'cricinfo.com', 'www.newindianexpress.com', 'www.nbmcw.com', 'timesofindia.indiatimes.com', 'www.newindianexpress.com', 'aircuttack.com', 'www.nbmcw.com', 'odishasuntimes.com', 'www.mapsofindia.com', 'www.sunhospitals.com', 'timesofindia.indiatimes.com', 'books.google.com', 'india9.com', 'books.google.com', 'www.nativeplanet.com', 'articles.economictimes.indiatimes.com', 'orissacinema.com', 'www.dailypioneer.com', 'baliyatra.org', 'www.srisriuniversity.org', 'www.svppgip.org', 'www.undp.org', 'www.odishastatemaritimemuseum.org', 'www.bpftio.org', 'www.osdma.org', ['2017 2nd international conference for convergence in technology ']]",1776398,Allow all users (no expiry set),101691,21 April 2005,202.62.226.149 ,2815,7,2005-04-21,2005-04,2005
666,666,Carmarthenshire,https://en.wikipedia.org/wiki/Carmarthenshire,51,2,"['10.2307/1790647', '10.1017/s0963926805002695', None, None, None, None]","[['the geographical journal'], ['urban history']]",3,5,0,20,0,0,21,0.058823529411764705,0.09803921568627451,0.39215686274509803,0.0392156862745098,0.0,0.19607843137254902,2,"['www.pembrokeshire.gov', 'legislation.gov', 'www.carmarthenshire.gov', 'www.carmarthenshire.gov', 'www.carmarthenshire.gov', 'www.abayoflife.com', 'books.google.com', 'www.discovercarmarthenshire.com', 'www.machynys.com', 'www.llansteffan.com', 'books.google.com', 'www.insidermedia.com', 'books.google.com', 'books.google.com', 'en.oxforddictionaries.com', 'www.abayoflife.com', 'books.google.com', 'www.penbontbren.com', 'www.discovercarmarthenshire.com', 'books.google.com', 'www.discovercarmarthenshire.com', 'primaryfacts.com', 'www.penbontbren.com', 'books.google.com', 'books.google.com', 'www.llandeilo.org', 'faw.org', 'histpop.org', ['the geographical journal'], ['urban history']]",154250,Allow all users (no expiry set),38669,4 December 2002,Renata ,618,1,2002-12-04,2002-12,2002
667,667,Legnano,https://en.wikipedia.org/wiki/Legnano,68,0,[],[],10,0,0,11,0,0,47,0.14705882352941177,0.0,0.16176470588235295,0.0,0.0,0.14705882352941177,0,"['cyclingranking.com', 'dolcegabbana.com', 'www.eurometeo.com', 'www.com', 'eurometeo.com', 'www.com', 'www.com', 'www.wunderground.com', 'sanmagno.com', 'www.com', 'www.legnanonews.com', 'consorziofiumeolona.org', 'legnano.org', 'legnano.org', 'earth-prints.org', 'legnano.org', 'legnano.org', 'legnano.org', 'www.legnano.org', 'legnano.org', 'legnano.org']",921430,Allow all users (no expiry set),97460,22 August 2004,ClockworkLunch ,481,0,2004-08-22,2004-08,2004
668,668,Cantabria,https://en.wikipedia.org/wiki/Cantabria,38,1,"['10.3989/aespa.085.012.008', None, None]",[['archivo español de arqueología']],3,0,0,7,0,0,27,0.07894736842105263,0.0,0.18421052631578946,0.02631578947368421,0.0,0.10526315789473684,1,"['www.etymonline.com', 'etymonline.com', 'www.etymonline.com', 'www.santandersummerfestival.com', 'www.collinsdictionary.com', 'www.ayto-selaya.com', 'www.festivalsantander.com', 'hdi.globaldatalab.org', 'es.wikisource.org', 'iso.org', ['archivo español de arqueología']]",69605,Allow all users (no expiry set),77885,9 August 2002,Perique des Palottes ,1348,1,2002-08-09,2002-08,2002
669,669,"Gubin, Poland","https://en.wikipedia.org/wiki/Gubin,_Poland",9,0,[],[],0,2,0,1,0,0,6,0.0,0.2222222222222222,0.1111111111111111,0.0,0.0,0.2222222222222222,0,"['www.gov', 'stat.gov', 'books.google.com']",703956,Allow all users (no expiry set),12579,4 June 2004,Cautious ,167,2,2004-06-04,2004-06,2004
670,670,Central Java,https://en.wikipedia.org/wiki/Central_Java,43,2,"['10.1126/science.7992059', '10.1146/annurev.an.17.100188.000355', '6410399', None, '384173', None]","[['periplus editions ltd ', 'annual review of anthropology ', 'proceedings of the national academy of sciences of the united states of america ', 'science magazine '], ['annual review of anthropology ']]",0,0,0,11,0,0,30,0.0,0.0,0.2558139534883721,0.046511627906976744,0.0,0.046511627906976744,2,"['wartakota.tribunnews.com', 'nasional.com', 'books.google.com', 'britannica.com', 'books.google.com', 'books.google.com', 'www.thejakartapost.com', 'www.kbri-bangkok.com', 'britannica.com', 'www.straitstimes.com', 'www.kompas.com', ['periplus editions ltd ', 'annual review of anthropology ', 'proceedings of the national academy of sciences of the united states of america ', 'science magazine '], ['annual review of anthropology ']]",453584,Allow all users (no expiry set),76768,3 February 2004,Morwen ,968,3,2004-02-03,2004-02,2004
671,671,Kalisz,https://en.wikipedia.org/wiki/Kalisz,40,3,"['10.1177/0265691417742017', '10.5194/hess-11-1633-2007', '10.1127/0941-2948/2006/0130', None, None, None, None, None, None]","[['european history quarterly'], ['hydrol. earth syst. sci. '], ['meteorologische zeitschrift']]",4,3,0,2,0,0,28,0.1,0.075,0.05,0.075,0.0,0.25,3,"['bdl.stat.gov', 'bdl.stat.gov', 'www.gov', 'www.google.com', 'www.google.com', 'encyclopedia.ushmm.org', 'yivoencyclopedia.org', 'encyclopedia.ushmm.org', 'sztetl.org', ['european history quarterly'], ['hydrol. earth syst. sci. '], ['meteorologische zeitschrift']]",74615,Allow all users (no expiry set),41568,22 August 2002,217.99.105.223 ,578,7,2002-08-22,2002-08,2002
672,672,Castel Goffredo,https://en.wikipedia.org/wiki/Castel_Goffredo,2,0,[],[],0,0,0,0,0,0,2,0.0,0.0,0.0,0.0,0.0,0.0,0,[],1050994,Allow all users (no expiry set),7899,8 October 2004,Pumpie ,125,0,2004-10-08,2004-10,2004
673,673,Bareq,https://en.wikipedia.org/wiki/Bareq,30,0,[],[],0,0,0,26,0,0,4,0.0,0.0,0.8666666666666667,0.0,0.0,0.0,0,"['books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.worldweatheronline.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com', 'books.google.com']",35582091,Allow all users (no expiry set),17706,22 April 2012,Zahiralbarqi ,295,0,2012-04-22,2012-04,2012
674,674,Capena,https://en.wikipedia.org/wiki/Capena,31,0,[],[],0,0,0,14,0,0,17,0.0,0.0,0.45161290322580644,0.0,0.0,0.0,0,"['olivecrona.wordpress.com', 'www.com', 'www.casacapena.com', 'blogs.laweekly.com', 'www.com', 'www.casacapena.com', 'www.travelpod.com', 'olivecrona.wordpress.com', 'www.com', 'www.capenaannozero.com', 'www.youtube.com', 'www.youtube.com', 'www.casacapena.com', 'www.com']",2687764,Allow all users (no expiry set),18808,16 September 2005,Water Bottle ,194,0,2005-09-16,2005-09,2005
675,675,Anabaptist–Jewish relations,https://en.wikipedia.org/wiki/Anabaptist%E2%80%93Jewish_relations,33,0,[],[],9,0,0,17,0,1,6,0.2727272727272727,0.0,0.5151515151515151,0.0,0.0,0.2727272727272727,0,"['www.etonline.com', 'forward.com', 'www.chicagotribune.com', 'www.mcall.com', 'www.nytimes.com', 'www.jpost.com', 'www.deseret.com', 'www.jpost.com', 'amishacres.com', 'www.vice.com', 'books.google.com', 'books.google.com', 'decentfilms.com', 'variety.com', 'www.jweekly.com', 'books.google.com', 'www.amazon.com', 'www.mennoworld.org', 'www.mennoworld.org', 'www.mennohof.org', 'www.yiddishbookcenter.org', 'oukosher.org', 'themennonite.org', 'sholemaleichem.org', 'www.splcenter.org', 'themennonite.org']",62110029,Allow all users (no expiry set),25661,20 October 2019,Bohemian Baltimore ,72,2,2019-10-20,2019-10,2019
676,676,Amasya,https://en.wikipedia.org/wiki/Amasya,24,1,[],[],2,1,0,5,0,0,15,0.08333333333333333,0.041666666666666664,0.20833333333333334,0.041666666666666664,0.0,0.16666666666666666,0,"['www.mgm.gov', 'books.google.com', 'jewishencyclopedia.com', 'www.hurriyetdailynews.com', 'books.google.com', 'books.google.com', 'www.catholic-hierarchy.org', 'cts.perseids.org']",1325621,Allow all users (no expiry set),48017,25 December 2004,OneGuy ,952,1,2004-12-25,2004-12,2004
677,677,Outline of Tunisia,https://en.wikipedia.org/wiki/Outline_of_Tunisia,1,0,[],[],0,1,0,0,0,0,0,0.0,1.0,0.0,0.0,0.0,1.0,0,['www.cia.gov'],16285795,Allow all users (no expiry set),22077,14 March 2008,The Transhumanist ,261,0,2008-03-14,2008-03,2008
678,678,Culture of Sussex,https://en.wikipedia.org/wiki/Culture_of_Sussex,142,1,[],[],26,4,0,21,0,6,84,0.18309859154929578,0.028169014084507043,0.14788732394366197,0.007042253521126761,0.0,0.21830985915492956,0,"['www.lewes.gov', 'www.southdowns.gov', 'www.eastsussex.gov', 'www.chichester.gov', 'www.bennettsassociates.com', 'www.britannica.com', 'www.thechampagnecompany.com', 'www.visitoruk.com', 'brightonfilm.com', 'www.cricinfo.com', 'historicalfoods.com', 'history-tourist.com', 'theculturetrip.com', 'historicalfoods.com', 'content.yudu.com', 'www.britainunlimited.com', 'findarticles.com', 'historicalfoods.com', 'britishairwaysi360.com', 'www.thakehamquaker.com', 'books.google.com', 'travel.nationalgeographic.com', 'www.ukrockfestivals.com', 'historicalfoods.com', 'www.francisfrith.com', 'www.charleston.org', 'econjwatch.org', 'www.sussexarch.org', 'www.nobelprize.org', 'www.visitsussex.org', 'www.biodiversitysussex.org', 'hastingspride.org', 'www.britishmuseum.org', 'www.nobelprize.org', 'www.filmcitybrighton.org', 'www.pbs.org', 'ukflagregistry.org', 'www.sussexrecordsociety.org', 'www.worthingdownlanders.org', 'www.englandschristianheritage.org', 'pallant.org', 'www.scfl.org', 'www.pallant.org', 'www.westdean.org', 'www.mybrightonandhove.org', 'brightonpermaculture.org', 'www.brightonphil.org', 'rth.org', 'www.nobelprize.org', 'www.fondation-fyssen.org', 'www.nobelprize.org']",38376685,Allow all users (no expiry set),77926,30 January 2013,Peetred ,301,2,2013-01-30,2013-01,2013
679,679,Kępno,https://en.wikipedia.org/wiki/K%C4%99pno,10,0,[],[],0,2,0,0,0,0,8,0.0,0.2,0.0,0.0,0.0,0.2,0,"['www.gov', 'pw.ipn.gov']",829399,Allow all users (no expiry set),11263,16 July 2004,PolishPoliticians ,122,1,2004-07-16,2004-07,2004
680,680,Mundaka,https://en.wikipedia.org/wiki/Mundaka,0,0,[],[],0,0,0,0,0,0,0,,,,,,,0,[],2883015,Allow all users (no expiry set),17281,11 October 2005,80.58.48.170 ,162,1,2005-10-11,2005-10,2005
681,681,Culture of Coimbatore,https://en.wikipedia.org/wiki/Culture_of_Coimbatore,29,0,[],[],1,0,0,23,0,0,5,0.034482758620689655,0.0,0.7931034482758621,0.0,0.0,0.034482758620689655,0,"['www.hinduonnet.com', 'books.google.com', 'www.hindu.com', 'articles.timesofindia.indiatimes.com', 'books.google.com', 'articles.timesofindia.indiatimes.com', 'www.thehindubusinessline.com', 'newindianexpress.com', 'www.hinduonnet.com', 'tamilinews.com', 'articles.timesofindia.indiatimes.com', 'tamil.samayam.com', 'maalaimalar.com', 'www.moneycontrol.com', 'www.maalaimalar.com', 'www.thecityvisit.com', 'economictimes.indiatimes.com', 'www.expressindia.com', 'books.google.com', 'books.google.com', 'www.hindu.com', 'www.thehindu.com', 'books.google.com', 'aicmeu.org']",46250566,Allow all users (no expiry set),16512,28 March 2015,Magentic Manifestations ,69,4,2015-03-28,2015-03,2015
682,682,Cairo Montenotte,https://en.wikipedia.org/wiki/Cairo_Montenotte,24,0,[],[],3,0,0,0,0,0,21,0.125,0.0,0.0,0.0,0.0,0.125,0,"['it.wikipedia.org', 'usrocchettese.altervista.org', 'it.wikipedia.org']",6570125,Allow all users (no expiry set),33380,20 August 2006,Eubot ,103,1,2006-08-20,2006-08,2006
683,683,Béni Abbès,https://en.wikipedia.org/wiki/B%C3%A9ni_Abb%C3%A8s,151,0,[],[],14,16,0,53,0,0,69,0.09271523178807947,0.10596026490066225,0.3509933774834437,0.0,0.0,0.1986754966887417,0,"['www.wilaya-bechar.gov', 'www.wilaya-bechar.gov', 'www.wilaya-bechar.gov', 'www.wilaya-bechar.gov', 'www.wilaya-bechar.gov', 'www.wilaya-bechar.gov', 'www.wilaya-bechar.gov', 'www.wilaya-bechar.gov', 'ftp.atdd.noaa.gov', 'www.wilaya-bechar.gov', 'www.wilaya-bechar.gov', 'www.wilaya-bechar.gov', 'www.wilaya-bechar.gov', 'www.wilaya-bechar.gov', 'www.wilaya-bechar.gov', 'www.wilaya-bechar.gov', 'books.google.com', 'www.saha-beniabbes.com', 'allocine.com', 'cache:nzgbu4uxg8ej:www.sonatrach-dz.com', 'www.algeriantourism.com', 'www.saha-beniabbes.com', 'www.mondomix.com', 'www.lesafriques.com', 'metz.consulat-algerie.com', 'saoura.over-blog.com', 'docs.google.com', 'saha-beniabbes.com', 'www.politiquemania.com', 'books.google.com', 'ayacom.jeeran.com', 'www.liberte-algerie.com', 'saoura.over-blog.com', 'el_maya.mondomix.com', 'www.vitaminedz.com', 'www.elmoudjahid.com', 'www.saha-beniabbes.com', 'www.1novembre54.com', 'www.statoids.com', 'www.djazairess.com', 'cache:b3i5b3cvd8sj:www.latribune-online.com', 'docs.google.com', 'www.maghress.com', 'ennaharonline.com', 'www.transactiondalgerie.com', 'www.annales.com', 'books.google.com', 'www.algeriepyrenees.com', 'books.google.com', 'www.francomix.com', 'www.artnet.com', 'www.babelouedstory.com', 'books.google.com', 'books.google.com', 'books.google.com', 'www.nomade-aventure.com', 'www.vitaminedz.com', 'books.google.com', 'voyage-algerie.com', 'docs.google.com', 'books.google.com', 'books.google.com', 'ouledziyad.jeeran.com', 'rouiba-ville.kazeo.com', 'sahara-nature.com', 'books.google.com', 'books.google.com', 'jsk1946.forumactif.com', 'books.google.com', 'consulatoran.ambafrance.org', 'www.nuits-metis.org', 'allies.alliance21.org', 'www03.us.archive.org', 'www.naturevivante.org', 'www.naturevivante.org', 'www.annales.org', 'www.rcd-algerie.org', 'fas.org', 'cache:i127wwzgghgj:amisdebeniabbes.org', 'www.cissan.org', 'benbadis.org', 'gouraya.org', 'www.nuits-metis.org']",15454653,Allow all users (no expiry set),86676,27 January 2008,Trabelsiismail ,398,0,2008-01-27,2008-01,2008
